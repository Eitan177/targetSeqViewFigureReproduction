HERE
3203
JJ
HH
Inside_Start:106466371 Inside_End:106466949 OutSide_Start:106467465 Oustide_End:106467732 chro:chr14 SVtype:2 sup:17 Avg_Span:704 sumProb:inf
Inside_Start:106466542 Inside_End:106466542 OutSide_Start:107074677 Oustide_End:107074677 chro:chr14 SVtype:2 sup:1 Avg_Span:608135 sumProb:inf
Inside_Start:106471245 Inside_End:106471245 OutSide_Start:107136716 Oustide_End:107136716 chro:chr14 SVtype:2 sup:2 Avg_Span:665471 sumProb:inf
Inside_Start:106478015 Inside_End:106478414 OutSide_Start:106805016 Oustide_End:106805556 chro:chr14 SVtype:2 sup:9 Avg_Span:327077 sumProb:inf
Inside_Start:106477946 Inside_End:106478176 OutSide_Start:106829613 Oustide_End:106829678 chro:chr14 SVtype:2 sup:24 Avg_Span:351582 sumProb:inf
Inside_Start:106634739 Inside_End:106634762 OutSide_Start:107137710 Oustide_End:107137857 chro:chr14 SVtype:2 sup:2 Avg_Span:503033 sumProb:inf
Inside_Start:106691328 Inside_End:106691599 OutSide_Start:107183244 Oustide_End:107183300 chro:chr14 SVtype:2 sup:51 Avg_Span:491782 sumProb:inf
Inside_Start:106785330 Inside_End:106785632 OutSide_Start:106810117 Oustide_End:106810537 chro:chr14 SVtype:2 sup:43 Avg_Span:24736 sumProb:inf
Inside_Start:106790778 Inside_End:106790890 OutSide_Start:107048552 Oustide_End:107048731 chro:chr14 SVtype:2 sup:25 Avg_Span:257704 sumProb:inf
Inside_Start:106798319 Inside_End:106798573 OutSide_Start:107106458 Oustide_End:107106532 chro:chr14 SVtype:2 sup:3 Avg_Span:308028 sumProb:inf
Inside_Start:106798536 Inside_End:106798540 OutSide_Start:106823154 Oustide_End:106823159 chro:chr14 SVtype:2 sup:8 Avg_Span:24618 sumProb:inf
Inside_Start:106805000 Inside_End:106805220 OutSide_Start:106829554 Oustide_End:106829646 chro:chr14 SVtype:2 sup:21 Avg_Span:24451 sumProb:inf
Inside_Start:106805114 Inside_End:106805222 OutSide_Start:106877523 Oustide_End:106877606 chro:chr14 SVtype:2 sup:27 Avg_Span:72421 sumProb:inf
Inside_Start:106804990 Inside_End:106805182 OutSide_Start:107094963 Oustide_End:107095212 chro:chr14 SVtype:2 sup:16 Avg_Span:290004 sumProb:inf
Inside_Start:106823078 Inside_End:106823082 OutSide_Start:107273698 Oustide_End:107273699 chro:chr14 SVtype:2 sup:4 Avg_Span:450618 sumProb:inf
Inside_Start:106993497 Inside_End:106993734 OutSide_Start:107183215 Oustide_End:107183307 chro:chr14 SVtype:2 sup:10 Avg_Span:189578 sumProb:inf
Inside_Start:107048497 Inside_End:107048650 OutSide_Start:107130926 Oustide_End:107131058 chro:chr14 SVtype:2 sup:14 Avg_Span:82398 sumProb:inf
Inside_Start:107057192 Inside_End:107057349 OutSide_Start:107275816 Oustide_End:107275861 chro:chr14 SVtype:2 sup:20 Avg_Span:218527 sumProb:inf
Inside_Start:32859651 Inside_End:32859673 OutSide_Start:33815661 Oustide_End:33815681 chro:chr16 SVtype:4 sup:2 Avg_Span:956009 sumProb:inf
Inside_Start:32993878 Inside_End:32994460 OutSide_Start:33673408 Oustide_End:33673699 chro:chr16 SVtype:4 sup:3 Avg_Span:679408 sumProb:inf
Inside_Start:97996616 Inside_End:97996754 OutSide_Start:98042142 Oustide_End:98042280 chro:chr2 SVtype:4 sup:2 Avg_Span:45526 sumProb:inf
Inside_Start:142493847 Inside_End:142494012 OutSide_Start:142510074 Oustide_End:142510173 chro:chr7 SVtype:4 sup:25 Avg_Span:16212 sumProb:25.000000
Inside_Start:22946661 Inside_End:22946733 OutSide_Start:22958493 Oustide_End:22958548 chro:chr14 SVtype:2 sup:16 Avg_Span:11813 sumProb:16.000000
Inside_Start:107239199 Inside_End:107239209 OutSide_Start:107239749 Oustide_End:107239924 chro:chr14 SVtype:2 sup:6 Avg_Span:647 sumProb:5.805264
Inside_Start:106653282 Inside_End:106653368 OutSide_Start:106845221 Oustide_End:106845297 chro:chr14 SVtype:2 sup:7 Avg_Span:191935 sumProb:4.998846
Inside_Start:106610194 Inside_End:106610307 OutSide_Start:106714307 Oustide_End:106714414 chro:chr14 SVtype:2 sup:5 Avg_Span:104110 sumProb:4.500000
Inside_Start:106674860 Inside_End:106674880 OutSide_Start:106933741 Oustide_End:106933788 chro:chr14 SVtype:2 sup:4 Avg_Span:258887 sumProb:4.000000
Inside_Start:106873470 Inside_End:106873470 OutSide_Start:106873878 Oustide_End:106873878 chro:chr14 SVtype:2 sup:4 Avg_Span:408 sumProb:4.000000
Inside_Start:107094868 Inside_End:107095014 OutSide_Start:107280866 Oustide_End:107280899 chro:chr14 SVtype:2 sup:26 Avg_Span:185946 sumProb:3.873658
Inside_Start:106477907 Inside_End:106478074 OutSide_Start:106780379 Oustide_End:106780596 chro:chr14 SVtype:2 sup:4 Avg_Span:302482 sumProb:3.264292
Inside_Start:106471005 Inside_End:106471032 OutSide_Start:107159672 Oustide_End:107159699 chro:chr14 SVtype:2 sup:3 Avg_Span:688658 sumProb:3.000000
Inside_Start:106518251 Inside_End:106518408 OutSide_Start:106573103 Oustide_End:106573287 chro:chr14 SVtype:2 sup:6 Avg_Span:54797 sumProb:3.000000
Inside_Start:106610223 Inside_End:106610278 OutSide_Start:107211005 Oustide_End:107211030 chro:chr14 SVtype:2 sup:3 Avg_Span:600760 sumProb:3.000000
Inside_Start:106669260 Inside_End:106669260 OutSide_Start:106928231 Oustide_End:106928231 chro:chr14 SVtype:2 sup:3 Avg_Span:258971 sumProb:3.000000
Inside_Start:106765104 Inside_End:106765104 OutSide_Start:106873830 Oustide_End:106873830 chro:chr14 SVtype:2 sup:3 Avg_Span:108726 sumProb:3.000000
Inside_Start:89161651 Inside_End:89161651 OutSide_Start:89197316 Oustide_End:89197316 chro:chr2 SVtype:5 sup:3 Avg_Span:35665 sumProb:3.000000
Inside_Start:142143360 Inside_End:142143360 OutSide_Start:142180232 Oustide_End:142180232 chro:chr7 SVtype:2 sup:3 Avg_Span:36872 sumProb:3.000000
Inside_Start:142138976 Inside_End:142139139 OutSide_Start:142157209 Oustide_End:142157238 chro:chr7 SVtype:2 sup:3 Avg_Span:18134 sumProb:2.999999
Inside_Start:106866125 Inside_End:106866417 OutSide_Start:107113616 Oustide_End:107113819 chro:chr14 SVtype:2 sup:4 Avg_Span:247459 sumProb:2.998802
Inside_Start:106518279 Inside_End:106518315 OutSide_Start:106725173 Oustide_End:106725236 chro:chr14 SVtype:2 sup:3 Avg_Span:206912 sumProb:2.997084
Inside_Start:106572947 Inside_End:106573210 OutSide_Start:106993619 Oustide_End:106993797 chro:chr14 SVtype:2 sup:4 Avg_Span:420632 sumProb:2.779514
Inside_Start:106350716 Inside_End:106350900 OutSide_Start:106360433 Oustide_End:106360533 chro:chr14 SVtype:2 sup:5 Avg_Span:9660 sumProb:2.387995
Inside_Start:89309479 Inside_End:89309529 OutSide_Start:89339764 Oustide_End:89339766 chro:chr2 SVtype:2 sup:3 Avg_Span:30253 sumProb:2.084691
Inside_Start:106873494 Inside_End:106873494 OutSide_Start:107148442 Oustide_End:107148442 chro:chr14 SVtype:2 sup:2 Avg_Span:274948 sumProb:2.021022
TOTAL 604
