HERE
3160
JJ
HH
Inside_Start:106478126 Inside_End:106478177 OutSide_Start:106780540 Oustide_End:106780562 chro:chr14 SVtype:2 sup:6 Avg_Span:302409 sumProb:inf
Inside_Start:106477882 Inside_End:106477958 OutSide_Start:107280990 Oustide_End:107281044 chro:chr14 SVtype:2 sup:3 Avg_Span:803109 sumProb:inf
Inside_Start:106518267 Inside_End:106518274 OutSide_Start:106691594 Oustide_End:106691609 chro:chr14 SVtype:2 sup:2 Avg_Span:173331 sumProb:inf
Inside_Start:106573036 Inside_End:106573300 OutSide_Start:107183318 Oustide_End:107183574 chro:chr14 SVtype:2 sup:7 Avg_Span:610276 sumProb:inf
Inside_Start:106573157 Inside_End:106573208 OutSide_Start:106691595 Oustide_End:106691723 chro:chr14 SVtype:2 sup:9 Avg_Span:118459 sumProb:inf
Inside_Start:106626902 Inside_End:106626902 OutSide_Start:107074681 Oustide_End:107074765 chro:chr14 SVtype:2 sup:2 Avg_Span:447821 sumProb:inf
Inside_Start:106691335 Inside_End:106691545 OutSide_Start:107183251 Oustide_End:107183302 chro:chr14 SVtype:2 sup:23 Avg_Span:491816 sumProb:inf
Inside_Start:106798311 Inside_End:106798539 OutSide_Start:106822930 Oustide_End:106823159 chro:chr14 SVtype:2 sup:4 Avg_Span:24619 sumProb:inf
Inside_Start:106798325 Inside_End:106798520 OutSide_Start:107106475 Oustide_End:107106504 chro:chr14 SVtype:2 sup:3 Avg_Span:308074 sumProb:inf
Inside_Start:106805108 Inside_End:106805225 OutSide_Start:107083057 Oustide_End:107083522 chro:chr14 SVtype:2 sup:27 Avg_Span:278114 sumProb:inf
Inside_Start:106805175 Inside_End:106805192 OutSide_Start:107095085 Oustide_End:107095273 chro:chr14 SVtype:2 sup:2 Avg_Span:289995 sumProb:inf
Inside_Start:106866162 Inside_End:106866445 OutSide_Start:107131018 Oustide_End:107131362 chro:chr14 SVtype:2 sup:10 Avg_Span:264775 sumProb:inf
Inside_Start:106993713 Inside_End:106993727 OutSide_Start:107183267 Oustide_End:107183315 chro:chr14 SVtype:2 sup:13 Avg_Span:189578 sumProb:inf
Inside_Start:107106246 Inside_End:107106411 OutSide_Start:107273699 Oustide_End:107273744 chro:chr14 SVtype:2 sup:3 Avg_Span:167410 sumProb:inf
Inside_Start:107148440 Inside_End:107148595 OutSide_Start:107169937 Oustide_End:107170173 chro:chr14 SVtype:2 sup:7 Avg_Span:21496 sumProb:inf
Inside_Start:32915350 Inside_End:32915350 OutSide_Start:33752304 Oustide_End:33752304 chro:chr16 SVtype:4 sup:4 Avg_Span:836954 sumProb:inf
Inside_Start:32990256 Inside_End:32990257 OutSide_Start:33677462 Oustide_End:33677462 chro:chr16 SVtype:4 sup:2 Avg_Span:687205 sumProb:inf
Inside_Start:32994110 Inside_End:32994459 OutSide_Start:33673410 Oustide_End:33673599 chro:chr16 SVtype:4 sup:8 Avg_Span:679153 sumProb:inf
Inside_Start:33021040 Inside_End:33021109 OutSide_Start:33647086 Oustide_End:33647152 chro:chr16 SVtype:4 sup:9 Avg_Span:626010 sumProb:inf
Inside_Start:32926975 Inside_End:32926981 OutSide_Start:33740687 Oustide_End:33740779 chro:chr16 SVtype:5 sup:2 Avg_Span:813755 sumProb:inf
Inside_Start:72004277 Inside_End:72004277 OutSide_Start:72156214 Oustide_End:72156214 chro:chrX SVtype:4 sup:2 Avg_Span:151937 sumProb:inf
Inside_Start:89442080 Inside_End:89442080 OutSide_Start:90078289 Oustide_End:90078289 chro:chr2 SVtype:4 sup:2 Avg_Span:636209 sumProb:inf
Inside_Start:89521086 Inside_End:89521197 OutSide_Start:89999544 Oustide_End:89999652 chro:chr2 SVtype:4 sup:2 Avg_Span:478456 sumProb:inf
Inside_Start:89533412 Inside_End:89533653 OutSide_Start:89976168 Oustide_End:89976399 chro:chr2 SVtype:4 sup:16 Avg_Span:442862 sumProb:inf
Inside_Start:92006403 Inside_End:92006498 OutSide_Start:92222329 Oustide_End:92222419 chro:chr2 SVtype:4 sup:4 Avg_Span:215969 sumProb:inf
Inside_Start:91679562 Inside_End:91679562 OutSide_Start:92222499 Oustide_End:92222499 chro:chr2 SVtype:5 sup:2 Avg_Span:542937 sumProb:inf
Inside_Start:142099472 Inside_End:142099486 OutSide_Start:142247276 Oustide_End:142247306 chro:chr7 SVtype:2 sup:3 Avg_Span:147814 sumProb:inf
Inside_Start:107218424 Inside_End:107218675 OutSide_Start:107253809 Oustide_End:107254020 chro:chr14 SVtype:2 sup:81 Avg_Span:35290 sumProb:81.000000
Inside_Start:107048460 Inside_End:107048681 OutSide_Start:107083254 Oustide_End:107083440 chro:chr14 SVtype:2 sup:104 Avg_Span:34716 sumProb:57.553123
Inside_Start:23004351 Inside_End:23004503 OutSide_Start:23564819 Oustide_End:23564949 chro:chr14 SVtype:4 sup:18 Avg_Span:560443 sumProb:18.000000
Inside_Start:106877352 Inside_End:106877620 OutSide_Start:107083173 Oustide_End:107083364 chro:chr14 SVtype:2 sup:41 Avg_Span:205763 sumProb:15.115394
Inside_Start:106466431 Inside_End:106466946 OutSide_Start:106467393 Oustide_End:106467683 chro:chr14 SVtype:2 sup:15 Avg_Span:665 sumProb:14.950645
Inside_Start:107239199 Inside_End:107239203 OutSide_Start:107239749 Oustide_End:107239994 chro:chr14 SVtype:2 sup:8 Avg_Span:706 sumProb:7.999977
Inside_Start:107136563 Inside_End:107136613 OutSide_Start:107169956 Oustide_End:107170135 chro:chr14 SVtype:2 sup:5 Avg_Span:33427 sumProb:4.999869
Inside_Start:22448286 Inside_End:22448412 OutSide_Start:22482773 Oustide_End:22483116 chro:chr15 SVtype:2 sup:4 Avg_Span:34562 sumProb:4.000000
Inside_Start:22465975 Inside_End:22466109 OutSide_Start:22482830 Oustide_End:22482935 chro:chr15 SVtype:2 sup:4 Avg_Span:16854 sumProb:3.999997
Inside_Start:89475660 Inside_End:89475805 OutSide_Start:90025343 Oustide_End:90025419 chro:chr2 SVtype:4 sup:11 Avg_Span:549642 sumProb:3.366225
Inside_Start:106825025 Inside_End:106825025 OutSide_Start:107022115 Oustide_End:107022115 chro:chr14 SVtype:2 sup:3 Avg_Span:197090 sumProb:3.000000
Inside_Start:107127639 Inside_End:107127653 OutSide_Start:107147909 Oustide_End:107148479 chro:chr14 SVtype:2 sup:3 Avg_Span:20645 sumProb:3.000000
Inside_Start:53724585 Inside_End:53724585 OutSide_Start:53724657 Oustide_End:53724657 chro:chr4 SVtype:5 sup:3 Avg_Span:72 sumProb:3.000000
Inside_Start:142028819 Inside_End:142028843 OutSide_Start:142161881 Oustide_End:142162110 chro:chr7 SVtype:5 sup:3 Avg_Span:133206 sumProb:3.000000
Inside_Start:142161618 Inside_End:142161895 OutSide_Start:142180241 Oustide_End:142180635 chro:chr7 SVtype:2 sup:3 Avg_Span:18701 sumProb:3.000000
Inside_Start:106597820 Inside_End:106597820 OutSide_Start:106798518 Oustide_End:106798518 chro:chr14 SVtype:2 sup:3 Avg_Span:200698 sumProb:2.999100
Inside_Start:2607558 Inside_End:2607558 OutSide_Start:2692640 Oustide_End:2692640 chro:chr16 SVtype:4 sup:3 Avg_Span:85082 sumProb:2.994643
Inside_Start:32859343 Inside_End:32859651 OutSide_Start:33815680 Oustide_End:33815730 chro:chr16 SVtype:4 sup:8 Avg_Span:956118 sumProb:2.724210
Inside_Start:107094790 Inside_End:107094999 OutSide_Start:107280872 Oustide_End:107280969 chro:chr14 SVtype:2 sup:15 Avg_Span:185957 sumProb:2.375993
Inside_Start:89609622 Inside_End:89609622 OutSide_Start:89891213 Oustide_End:89891213 chro:chr2 SVtype:4 sup:4 Avg_Span:281591 sumProb:2.297945
Inside_Start:106866091 Inside_End:106866399 OutSide_Start:107048539 Oustide_End:107048778 chro:chr14 SVtype:2 sup:38 Avg_Span:182316 sumProb:2.008604
Inside_Start:106653166 Inside_End:106653225 OutSide_Start:106866320 Oustide_End:106866330 chro:chr14 SVtype:2 sup:4 Avg_Span:213129 sumProb:2.000140
TOTAL 781
