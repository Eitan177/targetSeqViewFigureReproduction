HERE
2357
JJ
HH
Inside_Start:106466233 Inside_End:106466764 OutSide_Start:106467211 Oustide_End:106467753 chro:chr14 SVtype:2 sup:12 Avg_Span:562 sumProb:inf
Inside_Start:106477941 Inside_End:106478143 OutSide_Start:106829620 Oustide_End:106829683 chro:chr14 SVtype:2 sup:16 Avg_Span:351599 sumProb:inf
Inside_Start:106518103 Inside_End:106518449 OutSide_Start:106993610 Oustide_End:106993891 chro:chr14 SVtype:2 sup:9 Avg_Span:475477 sumProb:inf
Inside_Start:106785332 Inside_End:106785418 OutSide_Start:106810130 Oustide_End:106810532 chro:chr14 SVtype:2 sup:10 Avg_Span:24798 sumProb:inf
Inside_Start:106804998 Inside_End:106805175 OutSide_Start:106877530 Oustide_End:106877650 chro:chr14 SVtype:2 sup:15 Avg_Span:72467 sumProb:inf
Inside_Start:106804936 Inside_End:106805164 OutSide_Start:107083075 Oustide_End:107083401 chro:chr14 SVtype:2 sup:8 Avg_Span:278159 sumProb:inf
Inside_Start:107048334 Inside_End:107048559 OutSide_Start:107130899 Oustide_End:107131041 chro:chr14 SVtype:2 sup:3 Avg_Span:82519 sumProb:inf
Inside_Start:89160976 Inside_End:89160999 OutSide_Start:89197160 Oustide_End:89197213 chro:chr2 SVtype:4 sup:4 Avg_Span:36193 sumProb:inf
Inside_Start:142138944 Inside_End:142139141 OutSide_Start:142157195 Oustide_End:142157315 chro:chr7 SVtype:2 sup:7 Avg_Span:18179 sumProb:inf
Inside_Start:89161535 Inside_End:89161642 OutSide_Start:90078321 Oustide_End:90078398 chro:chr2 SVtype:5 sup:36 Avg_Span:916779 sumProb:21.701977
Inside_Start:106518043 Inside_End:106518227 OutSide_Start:107183231 Oustide_End:107183293 chro:chr14 SVtype:2 sup:21 Avg_Span:665070 sumProb:19.023882
Inside_Start:106691145 Inside_End:106691704 OutSide_Start:107183244 Oustide_End:107183435 chro:chr14 SVtype:2 sup:17 Avg_Span:491828 sumProb:17.009869
Inside_Start:107094858 Inside_End:107095064 OutSide_Start:107280870 Oustide_End:107281053 chro:chr14 SVtype:2 sup:18 Avg_Span:185963 sumProb:17.000034
Inside_Start:106993585 Inside_End:106993720 OutSide_Start:107183223 Oustide_End:107183337 chro:chr14 SVtype:2 sup:9 Avg_Span:189598 sumProb:9.022217
Inside_Start:106780296 Inside_End:106780451 OutSide_Start:107280878 Oustide_End:107281053 chro:chr14 SVtype:2 sup:12 Avg_Span:500596 sumProb:7.285240
Inside_Start:106572861 Inside_End:106572938 OutSide_Start:107183192 Oustide_End:107183301 chro:chr14 SVtype:2 sup:10 Avg_Span:610343 sumProb:7.068998
Inside_Start:23029836 Inside_End:23029944 OutSide_Start:23090502 Oustide_End:23091015 chro:chr22 SVtype:2 sup:7 Avg_Span:60812 sumProb:6.000003
Inside_Start:106866085 Inside_End:106866320 OutSide_Start:107048569 Oustide_End:107048609 chro:chr14 SVtype:2 sup:6 Avg_Span:182358 sumProb:5.993356
Inside_Start:106805003 Inside_End:106805061 OutSide_Start:107280947 Oustide_End:107280988 chro:chr14 SVtype:2 sup:5 Avg_Span:475929 sumProb:4.998802
Inside_Start:142143214 Inside_End:142143492 OutSide_Start:142180111 Oustide_End:142180502 chro:chr7 SVtype:2 sup:4 Avg_Span:36989 sumProb:4.000000
Inside_Start:106477827 Inside_End:106477942 OutSide_Start:107280918 Oustide_End:107280970 chro:chr14 SVtype:2 sup:4 Avg_Span:803057 sumProb:4.000000
Inside_Start:142111232 Inside_End:142111319 OutSide_Start:142131434 Oustide_End:142131569 chro:chr7 SVtype:2 sup:4 Avg_Span:20214 sumProb:3.998875
Inside_Start:33021099 Inside_End:33021133 OutSide_Start:33647059 Oustide_End:33647098 chro:chr16 SVtype:4 sup:4 Avg_Span:625979 sumProb:3.423074
Inside_Start:107083025 Inside_End:107083086 OutSide_Start:107280864 Oustide_End:107280928 chro:chr14 SVtype:2 sup:4 Avg_Span:197838 sumProb:3.291384
Inside_Start:106477865 Inside_End:106477903 OutSide_Start:106805133 Oustide_End:106805401 chro:chr14 SVtype:2 sup:3 Avg_Span:327370 sumProb:3.000003
Inside_Start:106626902 Inside_End:106627059 OutSide_Start:107074719 Oustide_End:107074820 chro:chr14 SVtype:2 sup:3 Avg_Span:447783 sumProb:3.000000
Inside_Start:107087240 Inside_End:107087269 OutSide_Start:107099220 Oustide_End:107099333 chro:chr14 SVtype:2 sup:4 Avg_Span:12007 sumProb:3.000000
Inside_Start:107122015 Inside_End:107122081 OutSide_Start:107198900 Oustide_End:107198984 chro:chr14 SVtype:2 sup:3 Avg_Span:76914 sumProb:3.000000
Inside_Start:142119736 Inside_End:142119860 OutSide_Start:142139263 Oustide_End:142139565 chro:chr7 SVtype:2 sup:3 Avg_Span:19615 sumProb:3.000000
Inside_Start:106653259 Inside_End:106653278 OutSide_Start:106845294 Oustide_End:106845339 chro:chr14 SVtype:2 sup:3 Avg_Span:192047 sumProb:2.997677
Inside_Start:32993849 Inside_End:32993901 OutSide_Start:33673674 Oustide_End:33673677 chro:chr16 SVtype:4 sup:3 Avg_Span:679809 sumProb:2.994870
Inside_Start:89399286 Inside_End:89399338 OutSide_Start:90193234 Oustide_End:90193272 chro:chr2 SVtype:4 sup:5 Avg_Span:793926 sumProb:2.989924
Inside_Start:106877620 Inside_End:106877692 OutSide_Start:107083285 Oustide_End:107083540 chro:chr14 SVtype:2 sup:5 Avg_Span:205785 sumProb:2.666960
Inside_Start:89619378 Inside_End:89619379 OutSide_Start:90121932 Oustide_End:90121938 chro:chr2 SVtype:4 sup:3 Avg_Span:502557 sumProb:2.486633
Inside_Start:106780309 Inside_End:106780372 OutSide_Start:107094984 Oustide_End:107095091 chro:chr14 SVtype:2 sup:3 Avg_Span:314669 sumProb:2.000525
Inside_Start:106518327 Inside_End:106518328 OutSide_Start:106573215 Oustide_End:106573216 chro:chr14 SVtype:2 sup:2 Avg_Span:54888 sumProb:2.000001
TOTAL 412
