HERE
12421
JJ
HH
Inside_Start:22997113 Inside_End:22997512 OutSide_Start:22997608 Oustide_End:22998024 chro:chr14 SVtype:2 sup:3 Avg_Span:478 sumProb:inf
Inside_Start:106466180 Inside_End:106466505 OutSide_Start:106466807 Oustide_End:106467543 chro:chr14 SVtype:2 sup:7 Avg_Span:888 sumProb:inf
Inside_Start:106466737 Inside_End:106467316 OutSide_Start:106467509 Oustide_End:106467910 chro:chr14 SVtype:2 sup:65 Avg_Span:681 sumProb:inf
Inside_Start:106477577 Inside_End:106478072 OutSide_Start:106780299 Oustide_End:106780939 chro:chr14 SVtype:2 sup:36 Avg_Span:302711 sumProb:inf
Inside_Start:106477695 Inside_End:106478067 OutSide_Start:106829589 Oustide_End:106829678 chro:chr14 SVtype:2 sup:23 Avg_Span:351666 sumProb:inf
Inside_Start:106691043 Inside_End:106691558 OutSide_Start:107183070 Oustide_End:107183608 chro:chr14 SVtype:2 sup:58 Avg_Span:491915 sumProb:inf
Inside_Start:106714261 Inside_End:106714302 OutSide_Start:106714685 Oustide_End:106714915 chro:chr14 SVtype:2 sup:2 Avg_Span:518 sumProb:inf
Inside_Start:106785021 Inside_End:106785517 OutSide_Start:106810114 Oustide_End:106810751 chro:chr14 SVtype:2 sup:52 Avg_Span:25002 sumProb:inf
Inside_Start:106797868 Inside_End:106798329 OutSide_Start:107106209 Oustide_End:107106735 chro:chr14 SVtype:2 sup:26 Avg_Span:308224 sumProb:inf
Inside_Start:106798031 Inside_End:106798630 OutSide_Start:106823158 Oustide_End:106823840 chro:chr14 SVtype:2 sup:96 Avg_Span:25117 sumProb:inf
Inside_Start:106804941 Inside_End:106805280 OutSide_Start:107083247 Oustide_End:107083759 chro:chr14 SVtype:2 sup:20 Avg_Span:278293 sumProb:inf
Inside_Start:106811299 Inside_End:106811801 OutSide_Start:106811822 Oustide_End:106812407 chro:chr14 SVtype:2 sup:31 Avg_Span:488 sumProb:inf
Inside_Start:106872910 Inside_End:106873336 OutSide_Start:106873349 Oustide_End:106873743 chro:chr14 SVtype:2 sup:10 Avg_Span:450 sumProb:inf
Inside_Start:107086636 Inside_End:107087230 OutSide_Start:107099002 Oustide_End:107099564 chro:chr14 SVtype:2 sup:21 Avg_Span:12153 sumProb:inf
Inside_Start:107087191 Inside_End:107087222 OutSide_Start:107113988 Oustide_End:107114005 chro:chr14 SVtype:2 sup:2 Avg_Span:26790 sumProb:inf
Inside_Start:107105940 Inside_End:107106391 OutSide_Start:107106398 Oustide_End:107106848 chro:chr14 SVtype:2 sup:12 Avg_Span:460 sumProb:inf
Inside_Start:22461204 Inside_End:22461763 OutSide_Start:22461777 Oustide_End:22462319 chro:chr15 SVtype:2 sup:11 Avg_Span:478 sumProb:inf
Inside_Start:32859007 Inside_End:32859607 OutSide_Start:33815129 Oustide_End:33815762 chro:chr16 SVtype:4 sup:40 Avg_Span:956225 sumProb:inf
Inside_Start:32994029 Inside_End:32994591 OutSide_Start:33672756 Oustide_End:33673408 chro:chr16 SVtype:4 sup:21 Avg_Span:678636 sumProb:inf
Inside_Start:31973269 Inside_End:31973867 OutSide_Start:32915259 Oustide_End:32915854 chro:chr16 SVtype:2 sup:29 Avg_Span:941924 sumProb:inf
Inside_Start:31974941 Inside_End:31975509 OutSide_Start:32916916 Oustide_End:32917422 chro:chr16 SVtype:2 sup:8 Avg_Span:941903 sumProb:inf
Inside_Start:31985799 Inside_End:31985854 OutSide_Start:32926864 Oustide_End:32926922 chro:chr16 SVtype:2 sup:7 Avg_Span:941066 sumProb:inf
Inside_Start:89495034 Inside_End:89495548 OutSide_Start:90025020 Oustide_End:90025594 chro:chr2 SVtype:4 sup:20 Avg_Span:529904 sumProb:inf
Inside_Start:89533098 Inside_End:89533685 OutSide_Start:89986441 Oustide_End:89987090 chro:chr2 SVtype:4 sup:34 Avg_Span:453393 sumProb:inf
Inside_Start:179954046 Inside_End:179954046 OutSide_Start:180467979 Oustide_End:180467979 chro:chr4 SVtype:2 sup:2 Avg_Span:513933 sumProb:inf
Inside_Start:1278190 Inside_End:1278755 OutSide_Start:1278778 Oustide_End:1279195 chro:chr5 SVtype:2 sup:12 Avg_Span:486 sumProb:inf
Inside_Start:106790401 Inside_End:106790922 OutSide_Start:106790925 Oustide_End:106791471 chro:chr14 SVtype:2 sup:106 Avg_Span:477 sumProb:49.120575
Inside_Start:106351303 Inside_End:106351733 OutSide_Start:106351740 Oustide_End:106352483 chro:chr14 SVtype:2 sup:37 Avg_Span:481 sumProb:36.994755
Inside_Start:107169454 Inside_End:107169950 OutSide_Start:107169963 Oustide_End:107170473 chro:chr14 SVtype:2 sup:36 Avg_Span:473 sumProb:36.217747
Inside_Start:107273434 Inside_End:107273870 OutSide_Start:107273870 Oustide_End:107274457 chro:chr14 SVtype:2 sup:34 Avg_Span:486 sumProb:33.999996
Inside_Start:106809931 Inside_End:106810374 OutSide_Start:106810378 Oustide_End:106810903 chro:chr14 SVtype:2 sup:34 Avg_Span:484 sumProb:33.000004
Inside_Start:106786721 Inside_End:106787272 OutSide_Start:106787274 Oustide_End:106787762 chro:chr14 SVtype:2 sup:33 Avg_Span:472 sumProb:30.498768
Inside_Start:107159404 Inside_End:107159893 OutSide_Start:107159899 Oustide_End:107160536 chro:chr14 SVtype:2 sup:30 Avg_Span:507 sumProb:29.999992
Inside_Start:33629727 Inside_End:33630191 OutSide_Start:33630194 Oustide_End:33630757 chro:chr16 SVtype:2 sup:30 Avg_Span:455 sumProb:28.999992
Inside_Start:89265137 Inside_End:89265668 OutSide_Start:89265672 Oustide_End:89266267 chro:chr2 SVtype:2 sup:29 Avg_Span:463 sumProb:28.250673
Inside_Start:89246382 Inside_End:89246802 OutSide_Start:89246872 Oustide_End:89247395 chro:chr2 SVtype:2 sup:32 Avg_Span:513 sumProb:27.484894
Inside_Start:22987164 Inside_End:22987696 OutSide_Start:22987709 Oustide_End:22988263 chro:chr14 SVtype:2 sup:27 Avg_Span:470 sumProb:27.000000
Inside_Start:106785208 Inside_End:106785689 OutSide_Start:106785713 Oustide_End:106786233 chro:chr14 SVtype:2 sup:32 Avg_Span:481 sumProb:26.410269
Inside_Start:106351750 Inside_End:106352239 OutSide_Start:106352248 Oustide_End:106352750 chro:chr14 SVtype:2 sup:26 Avg_Span:472 sumProb:26.049290
Inside_Start:106732613 Inside_End:106733122 OutSide_Start:106733128 Oustide_End:106733742 chro:chr14 SVtype:2 sup:26 Avg_Span:512 sumProb:26.000000
Inside_Start:106973900 Inside_End:106974375 OutSide_Start:106974384 Oustide_End:106975024 chro:chr14 SVtype:2 sup:26 Avg_Span:470 sumProb:26.000000
Inside_Start:106799620 Inside_End:106800185 OutSide_Start:106800198 Oustide_End:106800785 chro:chr14 SVtype:2 sup:32 Avg_Span:478 sumProb:25.287920
Inside_Start:22962212 Inside_End:22962714 OutSide_Start:22962727 Oustide_End:22963296 chro:chr14 SVtype:2 sup:25 Avg_Span:487 sumProb:25.000000
Inside_Start:22944752 Inside_End:22945287 OutSide_Start:22945294 Oustide_End:22945742 chro:chr14 SVtype:2 sup:24 Avg_Span:470 sumProb:24.000000
Inside_Start:22977559 Inside_End:22978073 OutSide_Start:22978073 Oustide_End:22978600 chro:chr14 SVtype:2 sup:23 Avg_Span:487 sumProb:23.000000
Inside_Start:107282407 Inside_End:107282891 OutSide_Start:107282916 Oustide_End:107283504 chro:chr14 SVtype:2 sup:23 Avg_Span:489 sumProb:22.997360
Inside_Start:22954514 Inside_End:22955020 OutSide_Start:22955044 Oustide_End:22955493 chro:chr14 SVtype:2 sup:22 Avg_Span:453 sumProb:22.000000
Inside_Start:22964392 Inside_End:22964898 OutSide_Start:22964916 Oustide_End:22965616 chro:chr14 SVtype:2 sup:22 Avg_Span:499 sumProb:22.000000
Inside_Start:22966196 Inside_End:22966603 OutSide_Start:22966677 Oustide_End:22967166 chro:chr14 SVtype:2 sup:22 Avg_Span:515 sumProb:22.000000
Inside_Start:23010583 Inside_End:23011041 OutSide_Start:23011100 Oustide_End:23011485 chro:chr14 SVtype:2 sup:22 Avg_Span:452 sumProb:22.000000
Inside_Start:23013436 Inside_End:23013892 OutSide_Start:23013906 Oustide_End:23014453 chro:chr14 SVtype:2 sup:22 Avg_Span:460 sumProb:22.000000
Inside_Start:106773581 Inside_End:106774013 OutSide_Start:106774044 Oustide_End:106774635 chro:chr14 SVtype:2 sup:22 Avg_Span:472 sumProb:22.000000
Inside_Start:106962582 Inside_End:106962930 OutSide_Start:106963016 Oustide_End:106963429 chro:chr14 SVtype:2 sup:22 Avg_Span:464 sumProb:22.000000
Inside_Start:107093042 Inside_End:107093358 OutSide_Start:107093635 Oustide_End:107093891 chro:chr14 SVtype:2 sup:22 Avg_Span:508 sumProb:22.000000
Inside_Start:106757179 Inside_End:106757593 OutSide_Start:106757599 Oustide_End:106758194 chro:chr14 SVtype:2 sup:22 Avg_Span:479 sumProb:21.999975
Inside_Start:107178217 Inside_End:107178744 OutSide_Start:107178824 Oustide_End:107179211 chro:chr14 SVtype:2 sup:22 Avg_Span:484 sumProb:21.998476
Inside_Start:89291355 Inside_End:89291809 OutSide_Start:89291815 Oustide_End:89292278 chro:chr2 SVtype:2 sup:29 Avg_Span:466 sumProb:21.492290
Inside_Start:106765015 Inside_End:106765580 OutSide_Start:106765586 Oustide_End:106766158 chro:chr14 SVtype:2 sup:21 Avg_Span:493 sumProb:21.000000
Inside_Start:106865822 Inside_End:106866329 OutSide_Start:106866343 Oustide_End:106866818 chro:chr14 SVtype:2 sup:21 Avg_Span:488 sumProb:20.989197
Inside_Start:23008477 Inside_End:23009001 OutSide_Start:23009016 Oustide_End:23009448 chro:chr14 SVtype:2 sup:20 Avg_Span:487 sumProb:20.000000
Inside_Start:107077969 Inside_End:107078405 OutSide_Start:107078426 Oustide_End:107079026 chro:chr14 SVtype:2 sup:20 Avg_Span:489 sumProb:20.000000
Inside_Start:107231429 Inside_End:107231844 OutSide_Start:107231892 Oustide_End:107232484 chro:chr14 SVtype:2 sup:20 Avg_Span:502 sumProb:20.000000
Inside_Start:22965195 Inside_End:22965621 OutSide_Start:22965742 Oustide_End:22966295 chro:chr14 SVtype:2 sup:20 Avg_Span:482 sumProb:19.998875
Inside_Start:91678784 Inside_End:91679350 OutSide_Start:91679353 Oustide_End:91679828 chro:chr2 SVtype:2 sup:122 Avg_Span:488 sumProb:19.536638
Inside_Start:20210744 Inside_End:20211323 OutSide_Start:20211323 Oustide_End:20211965 chro:chr15 SVtype:2 sup:69 Avg_Span:497 sumProb:19.092312
Inside_Start:106852027 Inside_End:106852455 OutSide_Start:106852458 Oustide_End:106852879 chro:chr14 SVtype:2 sup:19 Avg_Span:450 sumProb:19.000080
Inside_Start:106986326 Inside_End:106986800 OutSide_Start:106986800 Oustide_End:106987230 chro:chr14 SVtype:2 sup:19 Avg_Span:476 sumProb:19.000000
Inside_Start:107182733 Inside_End:107183178 OutSide_Start:107183203 Oustide_End:107183710 chro:chr14 SVtype:2 sup:19 Avg_Span:469 sumProb:18.990536
Inside_Start:22251289 Inside_End:22251666 OutSide_Start:22251731 Oustide_End:22252249 chro:chr14 SVtype:2 sup:18 Avg_Span:497 sumProb:18.000000
Inside_Start:106511169 Inside_End:106511622 OutSide_Start:106511658 Oustide_End:106512124 chro:chr14 SVtype:2 sup:18 Avg_Span:463 sumProb:18.000000
Inside_Start:107038829 Inside_End:107039302 OutSide_Start:107039334 Oustide_End:107039766 chro:chr14 SVtype:2 sup:18 Avg_Span:483 sumProb:18.000000
Inside_Start:107218069 Inside_End:107218598 OutSide_Start:107218610 Oustide_End:107219312 chro:chr14 SVtype:2 sup:19 Avg_Span:481 sumProb:17.999989
Inside_Start:106898563 Inside_End:106898989 OutSide_Start:106898992 Oustide_End:106899546 chro:chr14 SVtype:2 sup:18 Avg_Span:457 sumProb:17.994072
Inside_Start:106353715 Inside_End:106354134 OutSide_Start:106354169 Oustide_End:106354588 chro:chr14 SVtype:2 sup:18 Avg_Span:459 sumProb:17.925013
Inside_Start:107130398 Inside_End:107130963 OutSide_Start:107130973 Oustide_End:107131547 chro:chr14 SVtype:2 sup:22 Avg_Span:493 sumProb:17.489569
Inside_Start:89344958 Inside_End:89345507 OutSide_Start:90192752 Oustide_End:90193420 chro:chr2 SVtype:4 sup:46 Avg_Span:847822 sumProb:17.414078
Inside_Start:106780149 Inside_End:106780531 OutSide_Start:106780596 Oustide_End:106780977 chro:chr14 SVtype:2 sup:22 Avg_Span:460 sumProb:17.210344
Inside_Start:106350340 Inside_End:106350842 OutSide_Start:106350875 Oustide_End:106351274 chro:chr14 SVtype:2 sup:17 Avg_Span:453 sumProb:17.007732
Inside_Start:22986801 Inside_End:22987111 OutSide_Start:22987235 Oustide_End:22987565 chro:chr14 SVtype:2 sup:17 Avg_Span:458 sumProb:17.000000
Inside_Start:107055081 Inside_End:107055516 OutSide_Start:107055529 Oustide_End:107056026 chro:chr14 SVtype:2 sup:17 Avg_Span:464 sumProb:17.000000
Inside_Start:107147430 Inside_End:107147842 OutSide_Start:107147852 Oustide_End:107148295 chro:chr14 SVtype:2 sup:17 Avg_Span:452 sumProb:17.000000
Inside_Start:33605293 Inside_End:33605815 OutSide_Start:33605829 Oustide_End:33606251 chro:chr16 SVtype:2 sup:17 Avg_Span:446 sumProb:16.998863
Inside_Start:107056617 Inside_End:107057137 OutSide_Start:107057166 Oustide_End:107057613 chro:chr14 SVtype:2 sup:17 Avg_Span:486 sumProb:16.998035
Inside_Start:89596419 Inside_End:89597018 OutSide_Start:89923485 Oustide_End:89923997 chro:chr2 SVtype:4 sup:49 Avg_Span:327013 sumProb:16.229864
Inside_Start:22937591 Inside_End:22938004 OutSide_Start:22938004 Oustide_End:22938474 chro:chr14 SVtype:2 sup:16 Avg_Span:451 sumProb:16.000000
Inside_Start:22957055 Inside_End:22957638 OutSide_Start:22957706 Oustide_End:22958093 chro:chr14 SVtype:2 sup:16 Avg_Span:491 sumProb:16.000000
Inside_Start:22994093 Inside_End:22994547 OutSide_Start:22994562 Oustide_End:22995004 chro:chr14 SVtype:2 sup:16 Avg_Span:495 sumProb:16.000000
Inside_Start:106379859 Inside_End:106380359 OutSide_Start:106380365 Oustide_End:106380962 chro:chr14 SVtype:2 sup:16 Avg_Span:512 sumProb:16.000000
Inside_Start:22462152 Inside_End:22462565 OutSide_Start:22462632 Oustide_End:22463069 chro:chr15 SVtype:2 sup:16 Avg_Span:463 sumProb:16.000000
Inside_Start:107065342 Inside_End:107065770 OutSide_Start:107065806 Oustide_End:107066214 chro:chr14 SVtype:2 sup:16 Avg_Span:461 sumProb:15.998967
Inside_Start:106925675 Inside_End:106926110 OutSide_Start:106926117 Oustide_End:106926581 chro:chr14 SVtype:2 sup:16 Avg_Span:476 sumProb:15.998306
Inside_Start:89339108 Inside_End:89339705 OutSide_Start:90198652 Oustide_End:90199236 chro:chr2 SVtype:4 sup:38 Avg_Span:859480 sumProb:15.902744
Inside_Start:89629329 Inside_End:89629903 OutSide_Start:89890676 Oustide_End:89891310 chro:chr2 SVtype:4 sup:38 Avg_Span:261409 sumProb:15.540320
Inside_Start:89416233 Inside_End:89416816 OutSide_Start:90121556 Oustide_End:90122175 chro:chr2 SVtype:4 sup:52 Avg_Span:705269 sumProb:15.403172
Inside_Start:20212903 Inside_End:20213454 OutSide_Start:20213456 Oustide_End:20214060 chro:chr15 SVtype:2 sup:42 Avg_Span:478 sumProb:15.052418
Inside_Start:107041925 Inside_End:107042325 OutSide_Start:107042338 Oustide_End:107042794 chro:chr14 SVtype:2 sup:16 Avg_Span:478 sumProb:15.001408
Inside_Start:22508964 Inside_End:22509236 OutSide_Start:22509395 Oustide_End:22509715 chro:chr14 SVtype:2 sup:15 Avg_Span:450 sumProb:15.000010
Inside_Start:33618477 Inside_End:33618886 OutSide_Start:33618929 Oustide_End:33619466 chro:chr16 SVtype:2 sup:15 Avg_Span:496 sumProb:15.000009
Inside_Start:106944862 Inside_End:106945247 OutSide_Start:106945303 Oustide_End:106945772 chro:chr14 SVtype:2 sup:15 Avg_Span:450 sumProb:15.000000
Inside_Start:107280496 Inside_End:107280977 OutSide_Start:107280985 Oustide_End:107281465 chro:chr14 SVtype:2 sup:15 Avg_Span:459 sumProb:14.865482
Inside_Start:22969802 Inside_End:22970194 OutSide_Start:22970374 Oustide_End:22970648 chro:chr14 SVtype:2 sup:14 Avg_Span:497 sumProb:14.000000
Inside_Start:106372655 Inside_End:106373120 OutSide_Start:106373136 Oustide_End:106373625 chro:chr14 SVtype:2 sup:14 Avg_Span:479 sumProb:14.000000
Inside_Start:106873369 Inside_End:106873754 OutSide_Start:106873815 Oustide_End:106874269 chro:chr14 SVtype:2 sup:14 Avg_Span:477 sumProb:14.000000
Inside_Start:107112997 Inside_End:107113397 OutSide_Start:107113499 Oustide_End:107113863 chro:chr14 SVtype:2 sup:14 Avg_Span:477 sumProb:14.000000
Inside_Start:22465616 Inside_End:22466044 OutSide_Start:22466049 Oustide_End:22466580 chro:chr15 SVtype:2 sup:15 Avg_Span:465 sumProb:14.000000
Inside_Start:106378928 Inside_End:106379337 OutSide_Start:106379382 Oustide_End:106379773 chro:chr14 SVtype:2 sup:14 Avg_Span:461 sumProb:13.999989
Inside_Start:106370147 Inside_End:106370735 OutSide_Start:106370745 Oustide_End:106371249 chro:chr14 SVtype:2 sup:14 Avg_Span:484 sumProb:13.999985
Inside_Start:106652810 Inside_End:106653246 OutSide_Start:106653266 Oustide_End:106653730 chro:chr14 SVtype:2 sup:18 Avg_Span:471 sumProb:13.984344
Inside_Start:106798183 Inside_End:106798700 OutSide_Start:106798737 Oustide_End:106799156 chro:chr14 SVtype:2 sup:26 Avg_Span:530 sumProb:13.756436
Inside_Start:89567181 Inside_End:89567774 OutSide_Start:89952807 Oustide_End:89953421 chro:chr2 SVtype:4 sup:51 Avg_Span:385579 sumProb:13.509620
Inside_Start:20210332 Inside_End:20210783 OutSide_Start:20210788 Oustide_End:20211307 chro:chr15 SVtype:2 sup:41 Avg_Span:466 sumProb:13.354906
Inside_Start:21222786 Inside_End:21223187 OutSide_Start:21223200 Oustide_End:21223662 chro:chr15 SVtype:2 sup:35 Avg_Span:465 sumProb:13.354410
Inside_Start:22279676 Inside_End:22280106 OutSide_Start:22280200 Oustide_End:22280635 chro:chr14 SVtype:2 sup:13 Avg_Span:464 sumProb:13.000000
Inside_Start:22409438 Inside_End:22409866 OutSide_Start:22409876 Oustide_End:22410427 chro:chr14 SVtype:2 sup:13 Avg_Span:461 sumProb:13.000000
Inside_Start:22471430 Inside_End:22471732 OutSide_Start:22471904 Oustide_End:22472160 chro:chr14 SVtype:2 sup:13 Avg_Span:459 sumProb:13.000000
Inside_Start:22957705 Inside_End:22958278 OutSide_Start:22958345 Oustide_End:22958865 chro:chr14 SVtype:2 sup:13 Avg_Span:490 sumProb:13.000000
Inside_Start:22970832 Inside_End:22971201 OutSide_Start:22971243 Oustide_End:22971840 chro:chr14 SVtype:2 sup:13 Avg_Span:487 sumProb:13.000000
Inside_Start:22988545 Inside_End:22988956 OutSide_Start:22988967 Oustide_End:22989537 chro:chr14 SVtype:2 sup:13 Avg_Span:498 sumProb:13.000000
Inside_Start:23007263 Inside_End:23007678 OutSide_Start:23007764 Oustide_End:23008232 chro:chr14 SVtype:2 sup:13 Avg_Span:479 sumProb:13.000000
Inside_Start:33638002 Inside_End:33638486 OutSide_Start:33638498 Oustide_End:33639065 chro:chr9 SVtype:2 sup:13 Avg_Span:481 sumProb:13.000000
Inside_Start:106993449 Inside_End:106993815 OutSide_Start:106993896 Oustide_End:106994299 chro:chr14 SVtype:2 sup:14 Avg_Span:469 sumProb:12.992914
Inside_Start:106354196 Inside_End:106354668 OutSide_Start:106354675 Oustide_End:106355300 chro:chr14 SVtype:2 sup:13 Avg_Span:473 sumProb:12.986440
Inside_Start:89543639 Inside_End:89544208 OutSide_Start:89975995 Oustide_End:89976611 chro:chr2 SVtype:4 sup:37 Avg_Span:432417 sumProb:12.742846
Inside_Start:32077242 Inside_End:32077797 OutSide_Start:32077804 Oustide_End:32078451 chro:chr16 SVtype:2 sup:40 Avg_Span:495 sumProb:12.549355
Inside_Start:20208432 Inside_End:20208955 OutSide_Start:20208962 Oustide_End:20209478 chro:chr15 SVtype:2 sup:45 Avg_Span:456 sumProb:12.543974
Inside_Start:22974986 Inside_End:22975443 OutSide_Start:22975491 Oustide_End:22975996 chro:chr14 SVtype:2 sup:12 Avg_Span:497 sumProb:12.000070
Inside_Start:22111328 Inside_End:22111660 OutSide_Start:22111769 Oustide_End:22112125 chro:chr14 SVtype:2 sup:12 Avg_Span:437 sumProb:12.000000
Inside_Start:22433761 Inside_End:22434277 OutSide_Start:22434306 Oustide_End:22434732 chro:chr14 SVtype:2 sup:12 Avg_Span:482 sumProb:12.000000
Inside_Start:22446884 Inside_End:22447254 OutSide_Start:22447307 Oustide_End:22447735 chro:chr14 SVtype:2 sup:12 Avg_Span:464 sumProb:12.000000
Inside_Start:22616112 Inside_End:22616644 OutSide_Start:22616665 Oustide_End:22617147 chro:chr14 SVtype:2 sup:12 Avg_Span:479 sumProb:12.000000
Inside_Start:22962811 Inside_End:22963284 OutSide_Start:22963305 Oustide_End:22963820 chro:chr14 SVtype:2 sup:12 Avg_Span:512 sumProb:12.000000
Inside_Start:106346469 Inside_End:106347027 OutSide_Start:106347028 Oustide_End:106347511 chro:chr14 SVtype:2 sup:12 Avg_Span:457 sumProb:12.000000
Inside_Start:106832766 Inside_End:106833216 OutSide_Start:106833246 Oustide_End:106833755 chro:chr14 SVtype:2 sup:12 Avg_Span:483 sumProb:12.000000
Inside_Start:106966548 Inside_End:106967026 OutSide_Start:106967120 Oustide_End:106967504 chro:chr14 SVtype:2 sup:12 Avg_Span:486 sumProb:12.000000
Inside_Start:107107658 Inside_End:107108157 OutSide_Start:107108177 Oustide_End:107108696 chro:chr14 SVtype:2 sup:12 Avg_Span:489 sumProb:12.000000
Inside_Start:40745361 Inside_End:40745832 OutSide_Start:40745911 Oustide_End:40746287 chro:chr19 SVtype:2 sup:12 Avg_Span:465 sumProb:12.000000
Inside_Start:95629704 Inside_End:95630255 OutSide_Start:95630258 Oustide_End:95630841 chro:chr2 SVtype:2 sup:12 Avg_Span:472 sumProb:12.000000
Inside_Start:22320628 Inside_End:22321101 OutSide_Start:22321155 Oustide_End:22321604 chro:chr14 SVtype:2 sup:12 Avg_Span:461 sumProb:11.999998
Inside_Start:89308931 Inside_End:89309389 OutSide_Start:89309391 Oustide_End:89310138 chro:chr2 SVtype:2 sup:16 Avg_Span:471 sumProb:11.986586
Inside_Start:106551840 Inside_End:106552235 OutSide_Start:106552287 Oustide_End:106552785 chro:chr14 SVtype:2 sup:12 Avg_Span:475 sumProb:11.950954
Inside_Start:89618762 Inside_End:89619298 OutSide_Start:89901226 Oustide_End:89901917 chro:chr2 SVtype:4 sup:30 Avg_Span:282621 sumProb:11.917024
Inside_Start:107048279 Inside_End:107048550 OutSide_Start:107048686 Oustide_End:107049108 chro:chr14 SVtype:2 sup:13 Avg_Span:470 sumProb:11.483591
Inside_Start:89398873 Inside_End:89399365 OutSide_Start:89399370 Oustide_End:89399977 chro:chr2 SVtype:2 sup:19 Avg_Span:472 sumProb:11.126963
Inside_Start:21215711 Inside_End:21216305 OutSide_Start:21216311 Oustide_End:21216790 chro:chr15 SVtype:2 sup:34 Avg_Span:466 sumProb:11.087132
Inside_Start:22293595 Inside_End:22294062 OutSide_Start:22294187 Oustide_End:22294508 chro:chr14 SVtype:2 sup:11 Avg_Span:470 sumProb:11.000000
Inside_Start:22943708 Inside_End:22944105 OutSide_Start:22944154 Oustide_End:22944538 chro:chr14 SVtype:2 sup:11 Avg_Span:436 sumProb:11.000000
Inside_Start:22976422 Inside_End:22976676 OutSide_Start:22976842 Oustide_End:22977218 chro:chr14 SVtype:2 sup:11 Avg_Span:467 sumProb:11.000000
Inside_Start:106329033 Inside_End:106329529 OutSide_Start:106329558 Oustide_End:106330024 chro:chr14 SVtype:2 sup:11 Avg_Span:479 sumProb:11.000000
Inside_Start:106329959 Inside_End:106330511 OutSide_Start:106330525 Oustide_End:106330986 chro:chr14 SVtype:2 sup:11 Avg_Span:473 sumProb:11.000000
Inside_Start:106927788 Inside_End:106928172 OutSide_Start:106928216 Oustide_End:106928634 chro:chr14 SVtype:2 sup:11 Avg_Span:466 sumProb:11.000000
Inside_Start:107272996 Inside_End:107273369 OutSide_Start:107273443 Oustide_End:107273811 chro:chr14 SVtype:2 sup:11 Avg_Span:469 sumProb:11.000000
Inside_Start:33648980 Inside_End:33649548 OutSide_Start:33649648 Oustide_End:33650047 chro:chr9 SVtype:2 sup:11 Avg_Span:500 sumProb:11.000000
Inside_Start:33786452 Inside_End:33786953 OutSide_Start:33786958 Oustide_End:33787581 chro:chr9 SVtype:2 sup:11 Avg_Span:514 sumProb:11.000000
Inside_Start:106724488 Inside_End:106724942 OutSide_Start:106724946 Oustide_End:106725506 chro:chr14 SVtype:2 sup:11 Avg_Span:475 sumProb:10.999984
Inside_Start:33662138 Inside_End:33662517 OutSide_Start:33662731 Oustide_End:33663022 chro:chr9 SVtype:2 sup:11 Avg_Span:491 sumProb:10.999701
Inside_Start:106572610 Inside_End:106573134 OutSide_Start:106573139 Oustide_End:106573577 chro:chr14 SVtype:2 sup:13 Avg_Span:462 sumProb:10.998778
Inside_Start:106349019 Inside_End:106349612 OutSide_Start:106349643 Oustide_End:106350051 chro:chr14 SVtype:2 sup:12 Avg_Span:470 sumProb:10.853038
Inside_Start:107239200 Inside_End:107239634 OutSide_Start:107239845 Oustide_End:107240129 chro:chr14 SVtype:2 sup:11 Avg_Span:586 sumProb:10.133432
Inside_Start:98000298 Inside_End:98000868 OutSide_Start:98037486 Oustide_End:98038070 chro:chr2 SVtype:4 sup:25 Avg_Span:37137 sumProb:10.130829
Inside_Start:67047761 Inside_End:67048152 OutSide_Start:67048207 Oustide_End:67048572 chro:chr11 SVtype:2 sup:10 Avg_Span:449 sumProb:10.000000
Inside_Start:22392458 Inside_End:22392850 OutSide_Start:22392916 Oustide_End:22393390 chro:chr14 SVtype:2 sup:10 Avg_Span:464 sumProb:10.000000
Inside_Start:22675637 Inside_End:22676039 OutSide_Start:22676090 Oustide_End:22676524 chro:chr14 SVtype:2 sup:10 Avg_Span:480 sumProb:10.000000
Inside_Start:22694640 Inside_End:22695122 OutSide_Start:22695205 Oustide_End:22695640 chro:chr14 SVtype:2 sup:10 Avg_Span:480 sumProb:10.000000
Inside_Start:22946356 Inside_End:22946634 OutSide_Start:22946822 Oustide_End:22947046 chro:chr14 SVtype:2 sup:10 Avg_Span:453 sumProb:10.000000
Inside_Start:106330728 Inside_End:106331165 OutSide_Start:106331179 Oustide_End:106331681 chro:chr14 SVtype:2 sup:10 Avg_Span:480 sumProb:10.000000
Inside_Start:106331499 Inside_End:106331908 OutSide_Start:106331910 Oustide_End:106332346 chro:chr14 SVtype:2 sup:10 Avg_Span:442 sumProb:10.000000
Inside_Start:106369600 Inside_End:106370015 OutSide_Start:106370034 Oustide_End:106370463 chro:chr14 SVtype:2 sup:10 Avg_Span:465 sumProb:10.000000
Inside_Start:106880643 Inside_End:106881123 OutSide_Start:106881250 Oustide_End:106881572 chro:chr14 SVtype:2 sup:10 Avg_Span:471 sumProb:10.000000
Inside_Start:22460872 Inside_End:22461273 OutSide_Start:22461314 Oustide_End:22461736 chro:chr15 SVtype:2 sup:10 Avg_Span:449 sumProb:10.000000
Inside_Start:33682322 Inside_End:33682714 OutSide_Start:33682754 Oustide_End:33683237 chro:chr9 SVtype:2 sup:10 Avg_Span:479 sumProb:10.000000
Inside_Start:21216502 Inside_End:21216998 OutSide_Start:21217007 Oustide_End:21217453 chro:chr15 SVtype:2 sup:36 Avg_Span:448 sumProb:9.745438
Inside_Start:106811840 Inside_End:106812160 OutSide_Start:106812274 Oustide_End:106812679 chro:chr14 SVtype:2 sup:12 Avg_Span:490 sumProb:9.381823
Inside_Start:106377329 Inside_End:106377892 OutSide_Start:106377921 Oustide_End:106378323 chro:chr14 SVtype:2 sup:13 Avg_Span:472 sumProb:9.287758
Inside_Start:32908598 Inside_End:32909070 OutSide_Start:32909080 Oustide_End:32909552 chro:chr16 SVtype:2 sup:33 Avg_Span:486 sumProb:9.276430
Inside_Start:33020598 Inside_End:33021101 OutSide_Start:33646462 Oustide_End:33647098 chro:chr16 SVtype:4 sup:22 Avg_Span:625929 sumProb:9.129922
Inside_Start:22236743 Inside_End:22237168 OutSide_Start:22237326 Oustide_End:22237651 chro:chr14 SVtype:2 sup:9 Avg_Span:504 sumProb:9.000000
Inside_Start:22961888 Inside_End:22962210 OutSide_Start:22962324 Oustide_End:22962717 chro:chr14 SVtype:2 sup:9 Avg_Span:503 sumProb:9.000000
Inside_Start:23006010 Inside_End:23006446 OutSide_Start:23006467 Oustide_End:23006894 chro:chr14 SVtype:2 sup:9 Avg_Span:460 sumProb:9.000000
Inside_Start:106405157 Inside_End:106405537 OutSide_Start:106405584 Oustide_End:106405953 chro:chr14 SVtype:2 sup:9 Avg_Span:448 sumProb:9.000000
Inside_Start:106559219 Inside_End:106559538 OutSide_Start:106559686 Oustide_End:106560043 chro:chr14 SVtype:2 sup:9 Avg_Span:469 sumProb:9.000000
Inside_Start:107061810 Inside_End:107062098 OutSide_Start:107062220 Oustide_End:107062632 chro:chr14 SVtype:2 sup:9 Avg_Span:444 sumProb:9.000000
Inside_Start:107275435 Inside_End:107275815 OutSide_Start:107275926 Oustide_End:107276449 chro:chr14 SVtype:2 sup:9 Avg_Span:515 sumProb:9.000000
Inside_Start:90583637 Inside_End:90584146 OutSide_Start:90584147 Oustide_End:90584711 chro:chr9 SVtype:2 sup:9 Avg_Span:477 sumProb:9.000000
Inside_Start:106641037 Inside_End:106641528 OutSide_Start:106641532 Oustide_End:106642099 chro:chr14 SVtype:2 sup:10 Avg_Span:488 sumProb:8.999995
Inside_Start:107287239 Inside_End:107287609 OutSide_Start:107287645 Oustide_End:107288021 chro:chr14 SVtype:2 sup:9 Avg_Span:422 sumProb:8.999992
Inside_Start:106559377 Inside_End:106559528 OutSide_Start:107178808 Oustide_End:107179100 chro:chr14 SVtype:2 sup:9 Avg_Span:619463 sumProb:8.999659
Inside_Start:92005963 Inside_End:92006489 OutSide_Start:92221710 Oustide_End:92222340 chro:chr2 SVtype:4 sup:70 Avg_Span:215710 sumProb:8.836082
Inside_Start:106786582 Inside_End:106786773 OutSide_Start:106787118 Oustide_End:106787309 chro:chr14 SVtype:2 sup:9 Avg_Span:504 sumProb:8.821583
Inside_Start:107086878 Inside_End:107087443 OutSide_Start:107087445 Oustide_End:107087864 chro:chr14 SVtype:2 sup:13 Avg_Span:494 sumProb:8.499981
Inside_Start:89326202 Inside_End:89326657 OutSide_Start:89326719 Oustide_End:89327183 chro:chr2 SVtype:2 sup:14 Avg_Span:488 sumProb:8.372459
Inside_Start:106797862 Inside_End:106798162 OutSide_Start:106798387 Oustide_End:106798684 chro:chr14 SVtype:2 sup:21 Avg_Span:512 sumProb:8.359321
Inside_Start:89521070 Inside_End:89521572 OutSide_Start:89999668 Oustide_End:90000394 chro:chr2 SVtype:5 sup:35 Avg_Span:478570 sumProb:8.014851
Inside_Start:22192163 Inside_End:22192501 OutSide_Start:22192651 Oustide_End:22192949 chro:chr14 SVtype:2 sup:8 Avg_Span:481 sumProb:8.000000
Inside_Start:22386609 Inside_End:22387043 OutSide_Start:22387298 Oustide_End:22387571 chro:chr14 SVtype:2 sup:8 Avg_Span:521 sumProb:8.000000
Inside_Start:22539022 Inside_End:22539445 OutSide_Start:22539514 Oustide_End:22539921 chro:chr14 SVtype:2 sup:8 Avg_Span:482 sumProb:8.000000
Inside_Start:22591715 Inside_End:22592142 OutSide_Start:22592169 Oustide_End:22592587 chro:chr14 SVtype:2 sup:8 Avg_Span:445 sumProb:8.000000
Inside_Start:22689992 Inside_End:22690279 OutSide_Start:22690449 Oustide_End:22690744 chro:chr14 SVtype:2 sup:8 Avg_Span:472 sumProb:8.000000
Inside_Start:22771900 Inside_End:22772262 OutSide_Start:22772388 Oustide_End:22772833 chro:chr14 SVtype:2 sup:8 Avg_Span:529 sumProb:8.000000
Inside_Start:22978075 Inside_End:22978292 OutSide_Start:22978510 Oustide_End:22978761 chro:chr14 SVtype:2 sup:8 Avg_Span:440 sumProb:8.000000
Inside_Start:106379484 Inside_End:106379917 OutSide_Start:106379931 Oustide_End:106380325 chro:chr14 SVtype:2 sup:8 Avg_Span:446 sumProb:8.000000
Inside_Start:106501179 Inside_End:106501741 OutSide_Start:106501745 Oustide_End:106502197 chro:chr14 SVtype:2 sup:8 Avg_Span:496 sumProb:8.000000
Inside_Start:107127451 Inside_End:107127696 OutSide_Start:107127920 Oustide_End:107128156 chro:chr14 SVtype:2 sup:8 Avg_Span:486 sumProb:8.000000
Inside_Start:107258827 Inside_End:107259180 OutSide_Start:107259235 Oustide_End:107259616 chro:chr14 SVtype:2 sup:8 Avg_Span:436 sumProb:8.000000
Inside_Start:89160921 Inside_End:89161161 OutSide_Start:89161406 Oustide_End:89161587 chro:chr2 SVtype:2 sup:8 Avg_Span:477 sumProb:8.000000
Inside_Start:89185335 Inside_End:89185735 OutSide_Start:89185750 Oustide_End:89186201 chro:chr2 SVtype:2 sup:8 Avg_Span:461 sumProb:8.000000
Inside_Start:106347248 Inside_End:106347597 OutSide_Start:106347707 Oustide_End:106348063 chro:chr14 SVtype:2 sup:8 Avg_Span:458 sumProb:7.992650
Inside_Start:106652910 Inside_End:106653324 OutSide_Start:106845278 Oustide_End:106845702 chro:chr14 SVtype:2 sup:13 Avg_Span:192248 sumProb:7.976816
Inside_Start:97996201 Inside_End:97996732 OutSide_Start:98041579 Oustide_End:98042100 chro:chr2 SVtype:4 sup:33 Avg_Span:45413 sumProb:7.901993
Inside_Start:32993121 Inside_End:32993627 OutSide_Start:32993645 Oustide_End:32994184 chro:chr16 SVtype:2 sup:23 Avg_Span:479 sumProb:7.794106
Inside_Start:107074492 Inside_End:107074894 OutSide_Start:107074927 Oustide_End:107075349 chro:chr14 SVtype:2 sup:11 Avg_Span:467 sumProb:7.614725
Inside_Start:106804658 Inside_End:106805032 OutSide_Start:106805103 Oustide_End:106805635 chro:chr14 SVtype:2 sup:8 Avg_Span:509 sumProb:7.480027
Inside_Start:106691070 Inside_End:106691516 OutSide_Start:106691598 Oustide_End:106691934 chro:chr14 SVtype:2 sup:10 Avg_Span:460 sumProb:7.389509
Inside_Start:106368975 Inside_End:106369321 OutSide_Start:106369538 Oustide_End:106369780 chro:chr14 SVtype:2 sup:8 Avg_Span:517 sumProb:7.319625
Inside_Start:106790150 Inside_End:106790490 OutSide_Start:106790750 Oustide_End:106790914 chro:chr14 SVtype:2 sup:17 Avg_Span:469 sumProb:7.096629
Inside_Start:22090217 Inside_End:22090657 OutSide_Start:22090700 Oustide_End:22091094 chro:chr14 SVtype:2 sup:7 Avg_Span:465 sumProb:7.000000
Inside_Start:22337004 Inside_End:22337310 OutSide_Start:22337513 Oustide_End:22337794 chro:chr14 SVtype:2 sup:7 Avg_Span:487 sumProb:7.000000
Inside_Start:22356252 Inside_End:22356623 OutSide_Start:22356724 Oustide_End:22357277 chro:chr14 SVtype:2 sup:7 Avg_Span:502 sumProb:7.000000
Inside_Start:22475830 Inside_End:22476317 OutSide_Start:22476360 Oustide_End:22476769 chro:chr14 SVtype:2 sup:7 Avg_Span:504 sumProb:7.000000
Inside_Start:22520729 Inside_End:22521296 OutSide_Start:22521323 Oustide_End:22521707 chro:chr14 SVtype:2 sup:7 Avg_Span:490 sumProb:7.000000
Inside_Start:22580714 Inside_End:22581134 OutSide_Start:22581134 Oustide_End:22581707 chro:chr14 SVtype:2 sup:7 Avg_Span:473 sumProb:7.000000
Inside_Start:22733627 Inside_End:22733945 OutSide_Start:22734115 Oustide_End:22734382 chro:chr14 SVtype:2 sup:7 Avg_Span:478 sumProb:7.000000
Inside_Start:22944471 Inside_End:22944766 OutSide_Start:22945062 Oustide_End:22945214 chro:chr14 SVtype:2 sup:7 Avg_Span:474 sumProb:7.000000
Inside_Start:22947554 Inside_End:22947861 OutSide_Start:22948014 Oustide_End:22948340 chro:chr14 SVtype:2 sup:7 Avg_Span:486 sumProb:7.000000
Inside_Start:22984213 Inside_End:22984475 OutSide_Start:22984668 Oustide_End:22984993 chro:chr14 SVtype:2 sup:7 Avg_Span:458 sumProb:7.000000
Inside_Start:106493806 Inside_End:106494039 OutSide_Start:106494222 Oustide_End:106494541 chro:chr14 SVtype:2 sup:7 Avg_Span:470 sumProb:7.000000
Inside_Start:106602344 Inside_End:106602584 OutSide_Start:106602792 Oustide_End:106603048 chro:chr14 SVtype:2 sup:7 Avg_Span:445 sumProb:7.000000
Inside_Start:106986827 Inside_End:106987192 OutSide_Start:106987264 Oustide_End:106987756 chro:chr14 SVtype:2 sup:7 Avg_Span:500 sumProb:7.000000
Inside_Start:29994153 Inside_End:29994624 OutSide_Start:29994763 Oustide_End:29995092 chro:chr16 SVtype:2 sup:7 Avg_Span:466 sumProb:7.000000
Inside_Start:48113586 Inside_End:48114058 OutSide_Start:48114082 Oustide_End:48114518 chro:chr8 SVtype:2 sup:7 Avg_Span:513 sumProb:7.000000
Inside_Start:106346205 Inside_End:106346579 OutSide_Start:106346632 Oustide_End:106347003 chro:chr14 SVtype:2 sup:7 Avg_Span:452 sumProb:7.000000
Inside_Start:22988316 Inside_End:22988528 OutSide_Start:22988742 Oustide_End:22988936 chro:chr14 SVtype:2 sup:7 Avg_Span:430 sumProb:6.999995
Inside_Start:22465780 Inside_End:22466343 OutSide_Start:22466358 Oustide_End:22466750 chro:chr14 SVtype:2 sup:7 Avg_Span:487 sumProb:6.999887
Inside_Start:107034529 Inside_End:107034745 OutSide_Start:107034966 Oustide_End:107035177 chro:chr14 SVtype:2 sup:7 Avg_Span:447 sumProb:6.999358
Inside_Start:107198747 Inside_End:107198899 OutSide_Start:107199165 Oustide_End:107199378 chro:chr14 SVtype:2 sup:7 Avg_Span:441 sumProb:6.999264
Inside_Start:106350915 Inside_End:106351274 OutSide_Start:106351321 Oustide_End:106351850 chro:chr14 SVtype:2 sup:7 Avg_Span:493 sumProb:6.997422
Inside_Start:106666927 Inside_End:106667481 OutSide_Start:106667494 Oustide_End:106667898 chro:chr14 SVtype:2 sup:7 Avg_Span:475 sumProb:6.995020
Inside_Start:106349915 Inside_End:106350393 OutSide_Start:106350414 Oustide_End:106350827 chro:chr14 SVtype:2 sup:9 Avg_Span:463 sumProb:6.734294
Inside_Start:107082734 Inside_End:107083189 OutSide_Start:107083248 Oustide_End:107083598 chro:chr14 SVtype:2 sup:9 Avg_Span:453 sumProb:6.462051
Inside_Start:89384412 Inside_End:89384674 OutSide_Start:90153691 Oustide_End:90154006 chro:chr2 SVtype:4 sup:17 Avg_Span:769290 sumProb:6.327998
Inside_Start:89475150 Inside_End:89475731 OutSide_Start:90044005 Oustide_End:90044520 chro:chr2 SVtype:4 sup:35 Avg_Span:568909 sumProb:6.233435
Inside_Start:106375797 Inside_End:106376319 OutSide_Start:106376321 Oustide_End:106376723 chro:chr14 SVtype:2 sup:7 Avg_Span:466 sumProb:6.144410
Inside_Start:31973518 Inside_End:31973914 OutSide_Start:31973941 Oustide_End:31974430 chro:chr16 SVtype:2 sup:15 Avg_Span:504 sumProb:6.038082
Inside_Start:22180588 Inside_End:22180754 OutSide_Start:22181061 Oustide_End:22181167 chro:chr14 SVtype:2 sup:6 Avg_Span:432 sumProb:6.000000
Inside_Start:22740002 Inside_End:22740484 OutSide_Start:22740540 Oustide_End:22740952 chro:chr14 SVtype:2 sup:6 Avg_Span:486 sumProb:6.000000
Inside_Start:22958406 Inside_End:22958805 OutSide_Start:22958842 Oustide_End:22959236 chro:chr14 SVtype:2 sup:6 Avg_Span:473 sumProb:6.000000
Inside_Start:22995171 Inside_End:22995247 OutSide_Start:22995593 Oustide_End:22996068 chro:chr14 SVtype:2 sup:6 Avg_Span:539 sumProb:6.000000
Inside_Start:23012040 Inside_End:23012487 OutSide_Start:23012487 Oustide_End:23012948 chro:chr14 SVtype:2 sup:6 Avg_Span:442 sumProb:6.000000
Inside_Start:106375198 Inside_End:106375306 OutSide_Start:106375641 Oustide_End:106375832 chro:chr14 SVtype:2 sup:6 Avg_Span:463 sumProb:6.000000
Inside_Start:106538646 Inside_End:106539042 OutSide_Start:106539091 Oustide_End:106539464 chro:chr14 SVtype:2 sup:6 Avg_Span:441 sumProb:6.000000
Inside_Start:22482425 Inside_End:22482871 OutSide_Start:22482938 Oustide_End:22483341 chro:chr15 SVtype:2 sup:6 Avg_Span:472 sumProb:6.000000
Inside_Start:134885287 Inside_End:134885545 OutSide_Start:134885786 Oustide_End:134886013 chro:chr3 SVtype:2 sup:6 Avg_Span:491 sumProb:6.000000
Inside_Start:22965845 Inside_End:22966160 OutSide_Start:22966402 Oustide_End:22966573 chro:chr14 SVtype:2 sup:6 Avg_Span:488 sumProb:5.999999
Inside_Start:106331941 Inside_End:106332072 OutSide_Start:106332402 Oustide_End:106332604 chro:chr14 SVtype:2 sup:6 Avg_Span:459 sumProb:5.999998
Inside_Start:22447849 Inside_End:22448047 OutSide_Start:22448285 Oustide_End:22448497 chro:chr15 SVtype:2 sup:6 Avg_Span:456 sumProb:5.999995
Inside_Start:106828792 Inside_End:106829356 OutSide_Start:106829462 Oustide_End:106829871 chro:chr14 SVtype:2 sup:6 Avg_Span:495 sumProb:5.999967
Inside_Start:106804941 Inside_End:106805244 OutSide_Start:106877644 Oustide_End:106877661 chro:chr14 SVtype:2 sup:14 Avg_Span:72567 sumProb:5.950063
Inside_Start:33764171 Inside_End:33764542 OutSide_Start:33764623 Oustide_End:33765071 chro:chr16 SVtype:2 sup:12 Avg_Span:492 sumProb:5.543544
Inside_Start:21220186 Inside_End:21220643 OutSide_Start:21220678 Oustide_End:21221198 chro:chr15 SVtype:2 sup:21 Avg_Span:470 sumProb:5.482908
Inside_Start:106800228 Inside_End:106800464 OutSide_Start:106800690 Oustide_End:106800955 chro:chr14 SVtype:2 sup:11 Avg_Span:525 sumProb:5.466381
Inside_Start:106358889 Inside_End:106359288 OutSide_Start:106359332 Oustide_End:106359741 chro:chr14 SVtype:2 sup:8 Avg_Span:475 sumProb:5.375472
Inside_Start:23511757 Inside_End:23512241 OutSide_Start:23512249 Oustide_End:23512992 chro:chr15 SVtype:2 sup:19 Avg_Span:524 sumProb:5.306450
Inside_Start:22907673 Inside_End:22907910 OutSide_Start:22919078 Oustide_End:22919237 chro:chr14 SVtype:2 sup:5 Avg_Span:11344 sumProb:5.026784
Inside_Start:20216163 Inside_End:20216553 OutSide_Start:20216577 Oustide_End:20217094 chro:chr15 SVtype:2 sup:14 Avg_Span:479 sumProb:5.002421
Inside_Start:22554871 Inside_End:22555203 OutSide_Start:22555309 Oustide_End:22555739 chro:chr14 SVtype:2 sup:5 Avg_Span:486 sumProb:5.000000
Inside_Start:22631325 Inside_End:22631779 OutSide_Start:22631789 Oustide_End:22632198 chro:chr14 SVtype:2 sup:5 Avg_Span:449 sumProb:5.000000
Inside_Start:22927390 Inside_End:22927682 OutSide_Start:22927869 Oustide_End:22928163 chro:chr14 SVtype:2 sup:5 Avg_Span:479 sumProb:5.000000
Inside_Start:22963319 Inside_End:22963660 OutSide_Start:22963724 Oustide_End:22964172 chro:chr14 SVtype:2 sup:5 Avg_Span:536 sumProb:5.000000
Inside_Start:22976884 Inside_End:22977034 OutSide_Start:22977374 Oustide_End:22977498 chro:chr14 SVtype:2 sup:5 Avg_Span:470 sumProb:5.000000
Inside_Start:104751321 Inside_End:104751603 OutSide_Start:104751877 Oustide_End:104752123 chro:chr14 SVtype:2 sup:5 Avg_Span:516 sumProb:5.000000
Inside_Start:106329579 Inside_End:106329977 OutSide_Start:106329993 Oustide_End:106330422 chro:chr14 SVtype:2 sup:5 Avg_Span:432 sumProb:5.000000
Inside_Start:106356396 Inside_End:106356583 OutSide_Start:106356845 Oustide_End:106357064 chro:chr14 SVtype:2 sup:5 Avg_Span:457 sumProb:5.000000
Inside_Start:106384724 Inside_End:106385072 OutSide_Start:106385223 Oustide_End:106385656 chro:chr14 SVtype:2 sup:5 Avg_Span:475 sumProb:5.000000
Inside_Start:106470996 Inside_End:106471276 OutSide_Start:106471400 Oustide_End:106471688 chro:chr14 SVtype:2 sup:5 Avg_Span:441 sumProb:5.000000
Inside_Start:106668947 Inside_End:106669217 OutSide_Start:106669357 Oustide_End:106669702 chro:chr14 SVtype:2 sup:5 Avg_Span:453 sumProb:5.000000
Inside_Start:106751937 Inside_End:106752262 OutSide_Start:106752403 Oustide_End:106752732 chro:chr14 SVtype:2 sup:5 Avg_Span:460 sumProb:5.000000
Inside_Start:106774077 Inside_End:106774156 OutSide_Start:106774494 Oustide_End:106774638 chro:chr14 SVtype:2 sup:5 Avg_Span:454 sumProb:5.000000
Inside_Start:106852474 Inside_End:106852624 OutSide_Start:106852909 Oustide_End:106853077 chro:chr14 SVtype:2 sup:5 Avg_Span:432 sumProb:5.000000
Inside_Start:106877080 Inside_End:106877426 OutSide_Start:106877484 Oustide_End:106877919 chro:chr14 SVtype:2 sup:5 Avg_Span:449 sumProb:5.000000
Inside_Start:107146914 Inside_End:107147223 OutSide_Start:107147401 Oustide_End:107147699 chro:chr14 SVtype:2 sup:5 Avg_Span:470 sumProb:5.000000
Inside_Start:33629418 Inside_End:33629725 OutSide_Start:33629920 Oustide_End:33630177 chro:chr16 SVtype:2 sup:6 Avg_Span:493 sumProb:5.000000
Inside_Start:993651 Inside_End:994073 OutSide_Start:994096 Oustide_End:994496 chro:chr17 SVtype:2 sup:5 Avg_Span:456 sumProb:5.000000
Inside_Start:98017866 Inside_End:98018208 OutSide_Start:98018300 Oustide_End:98018702 chro:chr2 SVtype:2 sup:5 Avg_Span:443 sumProb:5.000000
Inside_Start:124520399 Inside_End:124520632 OutSide_Start:124520809 Oustide_End:124521049 chro:chr8 SVtype:2 sup:5 Avg_Span:444 sumProb:5.000000
Inside_Start:33629088 Inside_End:33629558 OutSide_Start:33629566 Oustide_End:33630004 chro:chr9 SVtype:2 sup:5 Avg_Span:446 sumProb:5.000000
Inside_Start:106382525 Inside_End:106382916 OutSide_Start:106382940 Oustide_End:106383380 chro:chr14 SVtype:2 sup:5 Avg_Span:446 sumProb:4.999987
Inside_Start:106724948 Inside_End:106725284 OutSide_Start:106725442 Oustide_End:106725856 chro:chr14 SVtype:2 sup:5 Avg_Span:472 sumProb:4.998875
Inside_Start:106381882 Inside_End:106382269 OutSide_Start:106382399 Oustide_End:106382781 chro:chr14 SVtype:2 sup:5 Avg_Span:483 sumProb:4.998865
Inside_Start:22964229 Inside_End:22964382 OutSide_Start:22964776 Oustide_End:22965054 chro:chr14 SVtype:2 sup:5 Avg_Span:545 sumProb:4.998045
Inside_Start:106993077 Inside_End:106993183 OutSide_Start:106993612 Oustide_End:106993839 chro:chr14 SVtype:2 sup:5 Avg_Span:557 sumProb:4.997308
Inside_Start:22372306 Inside_End:22372471 OutSide_Start:22372735 Oustide_End:22372956 chro:chr14 SVtype:2 sup:5 Avg_Span:470 sumProb:4.995345
Inside_Start:31963219 Inside_End:31963578 OutSide_Start:31963732 Oustide_End:31964053 chro:chr16 SVtype:2 sup:15 Avg_Span:475 sumProb:4.994823
Inside_Start:107150596 Inside_End:107150949 OutSide_Start:107151112 Oustide_End:107151429 chro:chr14 SVtype:2 sup:5 Avg_Span:480 sumProb:4.959966
Inside_Start:89512428 Inside_End:89512876 OutSide_Start:90007521 Oustide_End:90008262 chro:chr2 SVtype:4 sup:14 Avg_Span:495128 sumProb:4.839868
Inside_Start:95618493 Inside_End:95618901 OutSide_Start:95619007 Oustide_End:95619456 chro:chr2 SVtype:2 sup:5 Avg_Span:492 sumProb:4.831128
Inside_Start:32989720 Inside_End:32990296 OutSide_Start:33677067 Oustide_End:33677421 chro:chr16 SVtype:4 sup:36 Avg_Span:687401 sumProb:4.767715
Inside_Start:87565717 Inside_End:87566137 OutSide_Start:87566141 Oustide_End:87566576 chro:chr2 SVtype:2 sup:23 Avg_Span:461 sumProb:4.760062
Inside_Start:106518089 Inside_End:106518487 OutSide_Start:106518504 Oustide_End:106518924 chro:chr14 SVtype:2 sup:5 Avg_Span:447 sumProb:4.497803
Inside_Start:106865733 Inside_End:106866308 OutSide_Start:107048524 Oustide_End:107048601 chro:chr14 SVtype:2 sup:5 Avg_Span:182500 sumProb:4.088300
Inside_Start:106691294 Inside_End:106691480 OutSide_Start:106993609 Oustide_End:106993858 chro:chr14 SVtype:2 sup:4 Avg_Span:302300 sumProb:4.001749
Inside_Start:107174806 Inside_End:107175330 OutSide_Start:107175371 Oustide_End:107175823 chro:chr14 SVtype:2 sup:5 Avg_Span:486 sumProb:4.001012
Inside_Start:106898360 Inside_End:106898490 OutSide_Start:106898816 Oustide_End:106898917 chro:chr14 SVtype:2 sup:4 Avg_Span:472 sumProb:4.000000
Inside_Start:63698841 Inside_End:63698841 OutSide_Start:63701653 Oustide_End:63701653 chro:chr11 SVtype:2 sup:4 Avg_Span:2812 sumProb:4.000000
Inside_Start:69462463 Inside_End:69462811 OutSide_Start:69462880 Oustide_End:69463275 chro:chr11 SVtype:2 sup:4 Avg_Span:430 sumProb:4.000000
Inside_Start:108321134 Inside_End:108321582 OutSide_Start:108321630 Oustide_End:108322042 chro:chr12 SVtype:2 sup:4 Avg_Span:461 sumProb:4.000000
Inside_Start:22297742 Inside_End:22298138 OutSide_Start:22298209 Oustide_End:22298547 chro:chr14 SVtype:2 sup:4 Avg_Span:425 sumProb:4.000000
Inside_Start:22337599 Inside_End:22337717 OutSide_Start:22338088 Oustide_End:22338196 chro:chr14 SVtype:2 sup:4 Avg_Span:469 sumProb:4.000000
Inside_Start:22658583 Inside_End:22658837 OutSide_Start:22659024 Oustide_End:22659374 chro:chr14 SVtype:2 sup:4 Avg_Span:480 sumProb:4.000000
Inside_Start:22958898 Inside_End:22959057 OutSide_Start:22959382 Oustide_End:22959476 chro:chr14 SVtype:2 sup:4 Avg_Span:442 sumProb:4.000000
Inside_Start:22961229 Inside_End:22961472 OutSide_Start:22961639 Oustide_End:22961895 chro:chr14 SVtype:2 sup:4 Avg_Span:447 sumProb:4.000000
Inside_Start:103351526 Inside_End:103351807 OutSide_Start:103351958 Oustide_End:103352211 chro:chr14 SVtype:2 sup:4 Avg_Span:419 sumProb:4.000000
Inside_Start:106357273 Inside_End:106357445 OutSide_Start:106357751 Oustide_End:106357910 chro:chr14 SVtype:2 sup:4 Avg_Span:467 sumProb:4.000000
Inside_Start:106511664 Inside_End:106511826 OutSide_Start:106512070 Oustide_End:106512413 chro:chr14 SVtype:2 sup:4 Avg_Span:483 sumProb:4.000000
Inside_Start:106621292 Inside_End:106621576 OutSide_Start:106621733 Oustide_End:106622193 chro:chr14 SVtype:2 sup:5 Avg_Span:516 sumProb:4.000000
Inside_Start:106764990 Inside_End:106765108 OutSide_Start:106765444 Oustide_End:106765577 chro:chr14 SVtype:2 sup:4 Avg_Span:444 sumProb:4.000000
Inside_Start:106873849 Inside_End:106873892 OutSide_Start:106874283 Oustide_End:106874346 chro:chr14 SVtype:2 sup:4 Avg_Span:437 sumProb:4.000000
Inside_Start:107012380 Inside_End:107012514 OutSide_Start:107012784 Oustide_End:107012925 chro:chr14 SVtype:2 sup:4 Avg_Span:427 sumProb:4.000000
Inside_Start:107039418 Inside_End:107039501 OutSide_Start:107039909 Oustide_End:107039988 chro:chr14 SVtype:2 sup:4 Avg_Span:481 sumProb:4.000000
Inside_Start:107113621 Inside_End:107113774 OutSide_Start:107114074 Oustide_End:107114194 chro:chr14 SVtype:2 sup:4 Avg_Span:468 sumProb:4.000000
Inside_Start:107121979 Inside_End:107122110 OutSide_Start:107122480 Oustide_End:107122570 chro:chr14 SVtype:2 sup:4 Avg_Span:487 sumProb:4.000000
Inside_Start:107136517 Inside_End:107136645 OutSide_Start:107137001 Oustide_End:107137352 chro:chr14 SVtype:2 sup:4 Avg_Span:537 sumProb:4.000000
Inside_Start:107147869 Inside_End:107148219 OutSide_Start:107148293 Oustide_End:107148883 chro:chr14 SVtype:2 sup:4 Avg_Span:541 sumProb:4.000000
Inside_Start:33630202 Inside_End:33630299 OutSide_Start:33630656 Oustide_End:33630706 chro:chr16 SVtype:2 sup:4 Avg_Span:443 sumProb:4.000000
Inside_Start:11423723 Inside_End:11424092 OutSide_Start:11424136 Oustide_End:11424503 chro:chr1 SVtype:2 sup:4 Avg_Span:426 sumProb:4.000000
Inside_Start:33983183 Inside_End:33983514 OutSide_Start:33983648 Oustide_End:33983987 chro:chr1 SVtype:2 sup:4 Avg_Span:481 sumProb:4.000000
Inside_Start:104124210 Inside_End:104124624 OutSide_Start:104124821 Oustide_End:104125050 chro:chr8 SVtype:2 sup:4 Avg_Span:513 sumProb:4.000000
Inside_Start:33618025 Inside_End:33618199 OutSide_Start:33618553 Oustide_End:33618750 chro:chr9 SVtype:2 sup:4 Avg_Span:482 sumProb:4.000000
Inside_Start:107183208 Inside_End:107183303 OutSide_Start:107183647 Oustide_End:107183730 chro:chr14 SVtype:2 sup:4 Avg_Span:434 sumProb:3.999996
Inside_Start:106787360 Inside_End:106787787 OutSide_Start:106787795 Oustide_End:106788204 chro:chr14 SVtype:2 sup:5 Avg_Span:447 sumProb:3.999994
Inside_Start:106933353 Inside_End:106933778 OutSide_Start:107175334 Oustide_End:107175448 chro:chr14 SVtype:2 sup:5 Avg_Span:241781 sumProb:3.999993
Inside_Start:106824382 Inside_End:106824680 OutSide_Start:106824844 Oustide_End:106825110 chro:chr14 SVtype:2 sup:4 Avg_Span:436 sumProb:3.999993
Inside_Start:20226586 Inside_End:20226916 OutSide_Start:20227050 Oustide_End:20227358 chro:chr15 SVtype:2 sup:10 Avg_Span:468 sumProb:3.997279
Inside_Start:89459430 Inside_End:89459858 OutSide_Start:90060948 Oustide_End:90061519 chro:chr2 SVtype:5 sup:17 Avg_Span:601506 sumProb:3.962463
Inside_Start:89911315 Inside_End:89911677 OutSide_Start:89911779 Oustide_End:89912252 chro:chr2 SVtype:2 sup:13 Avg_Span:479 sumProb:3.925303
Inside_Start:89552352 Inside_End:89552947 OutSide_Start:89967241 Oustide_End:89967734 chro:chr2 SVtype:4 sup:9 Avg_Span:414790 sumProb:3.673854
Inside_Start:106378006 Inside_End:106378358 OutSide_Start:106378451 Oustide_End:106378892 chro:chr14 SVtype:2 sup:4 Avg_Span:461 sumProb:3.499580
Inside_Start:20270727 Inside_End:20271069 OutSide_Start:20271172 Oustide_End:20271866 chro:chr15 SVtype:2 sup:6 Avg_Span:615 sumProb:3.244352
Inside_Start:21217472 Inside_End:21217607 OutSide_Start:21217930 Oustide_End:21218087 chro:chr15 SVtype:2 sup:10 Avg_Span:449 sumProb:3.193234
Inside_Start:106790952 Inside_End:106791297 OutSide_Start:106816104 Oustide_End:106816514 chro:chr14 SVtype:2 sup:9 Avg_Span:25189 sumProb:3.190011
Inside_Start:32063081 Inside_End:32063669 OutSide_Start:33006766 Oustide_End:33007590 chro:chr16 SVtype:2 sup:20 Avg_Span:943720 sumProb:3.167363
Inside_Start:22489557 Inside_End:22489910 OutSide_Start:22490117 Oustide_End:22490464 chro:chr15 SVtype:2 sup:3 Avg_Span:556 sumProb:3.026138
Inside_Start:89629097 Inside_End:89629331 OutSide_Start:89891219 Oustide_End:89891367 chro:chr2 SVtype:4 sup:9 Avg_Span:262078 sumProb:3.016448
Inside_Start:89433995 Inside_End:89434491 OutSide_Start:90085340 Oustide_End:90085819 chro:chr2 SVtype:4 sup:7 Avg_Span:651219 sumProb:3.002665
Inside_Start:106465871 Inside_End:106466374 OutSide_Start:106467309 Oustide_End:106467550 chro:chr14 SVtype:2 sup:4 Avg_Span:1223 sumProb:3.002569
Inside_Start:21222483 Inside_End:21222655 OutSide_Start:21222944 Oustide_End:21223132 chro:chr15 SVtype:2 sup:10 Avg_Span:513 sumProb:3.000104
Inside_Start:106784942 Inside_End:106785004 OutSide_Start:106785536 Oustide_End:106785612 chro:chr14 SVtype:2 sup:3 Avg_Span:585 sumProb:3.000002
Inside_Start:106851837 Inside_End:106851937 OutSide_Start:106852351 Oustide_End:106852379 chro:chr14 SVtype:2 sup:3 Avg_Span:456 sumProb:3.000000
Inside_Start:127432352 Inside_End:127432352 OutSide_Start:127432798 Oustide_End:127432798 chro:chr10 SVtype:2 sup:3 Avg_Span:446 sumProb:3.000000
Inside_Start:60786475 Inside_End:60786875 OutSide_Start:60786985 Oustide_End:60787314 chro:chr11 SVtype:2 sup:3 Avg_Span:522 sumProb:3.000000
Inside_Start:64639032 Inside_End:64639289 OutSide_Start:64639468 Oustide_End:64639734 chro:chr11 SVtype:2 sup:3 Avg_Span:438 sumProb:3.000000
Inside_Start:67048280 Inside_End:67048302 OutSide_Start:67048695 Oustide_End:67048734 chro:chr11 SVtype:2 sup:3 Avg_Span:426 sumProb:3.000000
Inside_Start:100581749 Inside_End:100581982 OutSide_Start:100582300 Oustide_End:100582579 chro:chr12 SVtype:2 sup:3 Avg_Span:550 sumProb:3.000000
Inside_Start:125632448 Inside_End:125632867 OutSide_Start:125633009 Oustide_End:125633359 chro:chr12 SVtype:2 sup:3 Avg_Span:500 sumProb:3.000000
Inside_Start:53412938 Inside_End:53413252 OutSide_Start:53413400 Oustide_End:53413680 chro:chr13 SVtype:2 sup:3 Avg_Span:484 sumProb:3.000000
Inside_Start:22237461 Inside_End:22237508 OutSide_Start:22237867 Oustide_End:22238046 chro:chr14 SVtype:2 sup:3 Avg_Span:469 sumProb:3.000000
Inside_Start:22636483 Inside_End:22636645 OutSide_Start:22636957 Oustide_End:22637131 chro:chr14 SVtype:2 sup:3 Avg_Span:454 sumProb:3.000000
Inside_Start:22740627 Inside_End:22740637 OutSide_Start:22741063 Oustide_End:22741070 chro:chr14 SVtype:2 sup:3 Avg_Span:434 sumProb:3.000000
Inside_Start:22783227 Inside_End:22783609 OutSide_Start:22783890 Oustide_End:22784137 chro:chr14 SVtype:2 sup:3 Avg_Span:560 sumProb:3.000000
Inside_Start:22788891 Inside_End:22789095 OutSide_Start:22789481 Oustide_End:22789609 chro:chr14 SVtype:2 sup:3 Avg_Span:522 sumProb:3.000000
Inside_Start:22937466 Inside_End:22937550 OutSide_Start:22937896 Oustide_End:22937963 chro:chr14 SVtype:2 sup:3 Avg_Span:435 sumProb:3.000000
Inside_Start:22956120 Inside_End:22956186 OutSide_Start:22956661 Oustide_End:22956860 chro:chr14 SVtype:2 sup:3 Avg_Span:585 sumProb:3.000000
Inside_Start:22980948 Inside_End:22981394 OutSide_Start:22981568 Oustide_End:22981844 chro:chr14 SVtype:2 sup:3 Avg_Span:568 sumProb:3.000000
Inside_Start:22987714 Inside_End:22987769 OutSide_Start:22988179 Oustide_End:22988196 chro:chr14 SVtype:2 sup:3 Avg_Span:444 sumProb:3.000000
Inside_Start:22997735 Inside_End:22997998 OutSide_Start:22998194 Oustide_End:22998585 chro:chr14 SVtype:2 sup:3 Avg_Span:552 sumProb:3.000000
Inside_Start:23007890 Inside_End:23008051 OutSide_Start:23008328 Oustide_End:23008570 chro:chr14 SVtype:2 sup:3 Avg_Span:487 sumProb:3.000000
Inside_Start:23010462 Inside_End:23010529 OutSide_Start:23010905 Oustide_End:23011036 chro:chr14 SVtype:2 sup:3 Avg_Span:495 sumProb:3.000000
Inside_Start:23011117 Inside_End:23011150 OutSide_Start:23011537 Oustide_End:23011564 chro:chr14 SVtype:2 sup:3 Avg_Span:418 sumProb:3.000000
Inside_Start:106373275 Inside_End:106373343 OutSide_Start:106373691 Oustide_End:106373940 chro:chr14 SVtype:2 sup:3 Avg_Span:536 sumProb:3.000000
Inside_Start:106585572 Inside_End:106585984 OutSide_Start:106586143 Oustide_End:106586420 chro:chr14 SVtype:2 sup:3 Avg_Span:498 sumProb:3.000000
Inside_Start:106597556 Inside_End:106597828 OutSide_Start:106598015 Oustide_End:106598271 chro:chr14 SVtype:2 sup:3 Avg_Span:444 sumProb:3.000000
Inside_Start:106674570 Inside_End:106674879 OutSide_Start:106675020 Oustide_End:106675294 chro:chr14 SVtype:2 sup:3 Avg_Span:453 sumProb:3.000000
Inside_Start:106877507 Inside_End:106877917 OutSide_Start:106877970 Oustide_End:106878386 chro:chr14 SVtype:2 sup:3 Avg_Span:466 sumProb:3.000000
Inside_Start:106974388 Inside_End:106974473 OutSide_Start:106974853 Oustide_End:106974931 chro:chr14 SVtype:2 sup:3 Avg_Span:457 sumProb:3.000000
Inside_Start:106986085 Inside_End:106986284 OutSide_Start:106986528 Oustide_End:106986727 chro:chr14 SVtype:2 sup:3 Avg_Span:474 sumProb:3.000000
Inside_Start:107021975 Inside_End:107022035 OutSide_Start:107022388 Oustide_End:107022542 chro:chr14 SVtype:2 sup:3 Avg_Span:447 sumProb:3.000000
Inside_Start:107210818 Inside_End:107211093 OutSide_Start:107211254 Oustide_End:107211557 chro:chr14 SVtype:2 sup:3 Avg_Span:485 sumProb:3.000000
Inside_Start:107282921 Inside_End:107283517 OutSide_Start:107283519 Oustide_End:107283939 chro:chr14 SVtype:2 sup:3 Avg_Span:539 sumProb:3.000000
Inside_Start:22472888 Inside_End:22472960 OutSide_Start:22473363 Oustide_End:22473385 chro:chr15 SVtype:2 sup:3 Avg_Span:448 sumProb:3.000000
Inside_Start:28108122 Inside_End:28108122 OutSide_Start:28108559 Oustide_End:28108603 chro:chr15 SVtype:2 sup:3 Avg_Span:466 sumProb:3.000000
Inside_Start:29994814 Inside_End:29994960 OutSide_Start:29995284 Oustide_End:29995435 chro:chr16 SVtype:2 sup:3 Avg_Span:458 sumProb:3.000000
Inside_Start:11395789 Inside_End:11395950 OutSide_Start:11396263 Oustide_End:11396380 chro:chr17 SVtype:2 sup:3 Avg_Span:444 sumProb:3.000000
Inside_Start:41013384 Inside_End:41013720 OutSide_Start:41013829 Oustide_End:41014207 chro:chr17 SVtype:2 sup:3 Avg_Span:472 sumProb:3.000000
Inside_Start:76720554 Inside_End:76720952 OutSide_Start:76721144 Oustide_End:76721371 chro:chr17 SVtype:2 sup:3 Avg_Span:533 sumProb:3.000000
Inside_Start:80366776 Inside_End:80366961 OutSide_Start:80367215 Oustide_End:80367370 chro:chr17 SVtype:2 sup:3 Avg_Span:419 sumProb:3.000000
Inside_Start:9962778 Inside_End:9962923 OutSide_Start:9963316 Oustide_End:9963433 chro:chr19 SVtype:2 sup:3 Avg_Span:519 sumProb:3.000000
Inside_Start:40745997 Inside_End:40746019 OutSide_Start:40746441 Oustide_End:40746444 chro:chr19 SVtype:2 sup:3 Avg_Span:430 sumProb:3.000000
Inside_Start:61032999 Inside_End:61033352 OutSide_Start:61033513 Oustide_End:61033760 chro:chr20 SVtype:2 sup:3 Avg_Span:443 sumProb:3.000000
Inside_Start:95639536 Inside_End:95639744 OutSide_Start:95639972 Oustide_End:95640167 chro:chr2 SVtype:2 sup:3 Avg_Span:427 sumProb:3.000000
Inside_Start:134514258 Inside_End:134514440 OutSide_Start:134514724 Oustide_End:134514876 chro:chr3 SVtype:2 sup:3 Avg_Span:450 sumProb:3.000000
Inside_Start:197400114 Inside_End:197400114 OutSide_Start:197400590 Oustide_End:197400590 chro:chr3 SVtype:2 sup:3 Avg_Span:476 sumProb:3.000000
Inside_Start:38327706 Inside_End:38327897 OutSide_Start:38328139 Oustide_End:38328508 chro:chr4 SVtype:2 sup:3 Avg_Span:483 sumProb:3.000000
Inside_Start:190100269 Inside_End:190100269 OutSide_Start:190100683 Oustide_End:190100683 chro:chr4 SVtype:2 sup:3 Avg_Span:414 sumProb:3.000000
Inside_Start:679379 Inside_End:679379 OutSide_Start:771534 Oustide_End:771534 chro:chr5 SVtype:2 sup:3 Avg_Span:92155 sumProb:3.000000
Inside_Start:132017830 Inside_End:132018054 OutSide_Start:132018434 Oustide_End:132018537 chro:chr8 SVtype:2 sup:3 Avg_Span:563 sumProb:3.000000
Inside_Start:33695775 Inside_End:33695987 OutSide_Start:33696254 Oustide_End:33696555 chro:chr9 SVtype:2 sup:3 Avg_Span:502 sumProb:3.000000
Inside_Start:106573155 Inside_End:106573578 OutSide_Start:106573632 Oustide_End:106574034 chro:chr14 SVtype:2 sup:3 Avg_Span:469 sumProb:3.000000
Inside_Start:106866436 Inside_End:106866445 OutSide_Start:106866919 Oustide_End:106866963 chro:chr14 SVtype:2 sup:3 Avg_Span:499 sumProb:3.000000
Inside_Start:106626870 Inside_End:106627323 OutSide_Start:106627328 Oustide_End:106627797 chro:chr14 SVtype:2 sup:3 Avg_Span:472 sumProb:2.999999
Inside_Start:106517793 Inside_End:106517880 OutSide_Start:106518211 Oustide_End:106518290 chro:chr14 SVtype:2 sup:3 Avg_Span:425 sumProb:2.999999
Inside_Start:106372239 Inside_End:106372481 OutSide_Start:106372874 Oustide_End:106372940 chro:chr14 SVtype:2 sup:3 Avg_Span:523 sumProb:2.999999
Inside_Start:106844646 Inside_End:106844811 OutSide_Start:106845121 Oustide_End:106845286 chro:chr14 SVtype:2 sup:4 Avg_Span:493 sumProb:2.999998
Inside_Start:22982261 Inside_End:22982805 OutSide_Start:22982903 Oustide_End:22983245 chro:chr14 SVtype:2 sup:3 Avg_Span:511 sumProb:2.999948
Inside_Start:106865589 Inside_End:106865819 OutSide_Start:106866141 Oustide_End:106866314 chro:chr14 SVtype:2 sup:4 Avg_Span:480 sumProb:2.998685
Inside_Start:106370796 Inside_End:106370855 OutSide_Start:106371290 Oustide_End:106371506 chro:chr14 SVtype:2 sup:3 Avg_Span:543 sumProb:2.996749
Inside_Start:106733178 Inside_End:106733178 OutSide_Start:107048743 Oustide_End:107048743 chro:chr14 SVtype:2 sup:3 Avg_Span:315565 sumProb:2.995937
Inside_Start:106466393 Inside_End:106466420 OutSide_Start:106466827 Oustide_End:106466830 chro:chr14 SVtype:2 sup:3 Avg_Span:426 sumProb:2.975296
Inside_Start:42680600 Inside_End:42681163 OutSide_Start:42681177 Oustide_End:42681606 chro:chr10 SVtype:2 sup:8 Avg_Span:516 sumProb:2.799768
Inside_Start:20208982 Inside_End:20209133 OutSide_Start:20209405 Oustide_End:20209612 chro:chr15 SVtype:2 sup:8 Avg_Span:471 sumProb:2.750412
Inside_Start:33647220 Inside_End:33647469 OutSide_Start:33647683 Oustide_End:33647986 chro:chr16 SVtype:2 sup:9 Avg_Span:477 sumProb:2.744634
Inside_Start:106359511 Inside_End:106359859 OutSide_Start:106359932 Oustide_End:106360381 chro:chr14 SVtype:2 sup:3 Avg_Span:484 sumProb:2.612761
Inside_Start:89291505 Inside_End:89291871 OutSide_Start:90259626 Oustide_End:90260079 chro:chr2 SVtype:4 sup:9 Avg_Span:968195 sumProb:2.502522
Inside_Start:106799419 Inside_End:106799706 OutSide_Start:106799826 Oustide_End:106800128 chro:chr14 SVtype:2 sup:3 Avg_Span:426 sumProb:2.499996
Inside_Start:106815262 Inside_End:106815660 OutSide_Start:106815684 Oustide_End:106816134 chro:chr14 SVtype:2 sup:3 Avg_Span:440 sumProb:2.496173
Inside_Start:89953261 Inside_End:89953584 OutSide_Start:89953947 Oustide_End:89954190 chro:chr2 SVtype:2 sup:8 Avg_Span:589 sumProb:2.494602
Inside_Start:106477440 Inside_End:106477988 OutSide_Start:106478014 Oustide_End:106478437 chro:chr14 SVtype:2 sup:4 Avg_Span:513 sumProb:2.493944
Inside_Start:21218067 Inside_End:21218159 OutSide_Start:21218496 Oustide_End:21218754 chro:chr15 SVtype:2 sup:9 Avg_Span:468 sumProb:2.491715
Inside_Start:91679358 Inside_End:91679630 OutSide_Start:91679796 Oustide_End:91680076 chro:chr2 SVtype:2 sup:15 Avg_Span:454 sumProb:2.253364
Inside_Start:32050625 Inside_End:32051048 OutSide_Start:32051287 Oustide_End:32051478 chro:chr16 SVtype:2 sup:6 Avg_Span:500 sumProb:2.153227
Inside_Start:51864179 Inside_End:51864179 OutSide_Start:51864662 Oustide_End:51864662 chro:chr16 SVtype:2 sup:2 Avg_Span:483 sumProb:2.063540
Inside_Start:107148442 Inside_End:107148736 OutSide_Start:107148876 Oustide_End:107149150 chro:chr14 SVtype:2 sup:3 Avg_Span:420 sumProb:2.000761
Inside_Start:97716551 Inside_End:97716985 OutSide_Start:97717027 Oustide_End:97717397 chro:chr2 SVtype:2 sup:5 Avg_Span:450 sumProb:2.000589
Inside_Start:106477642 Inside_End:106478094 OutSide_Start:106877367 Oustide_End:106877655 chro:chr14 SVtype:2 sup:3 Avg_Span:399670 sumProb:2.000096
Inside_Start:107178878 Inside_End:107178888 OutSide_Start:107179459 Oustide_End:107179487 chro:chr14 SVtype:2 sup:2 Avg_Span:590 sumProb:2.000003
Inside_Start:74455301 Inside_End:74455301 OutSide_Start:74455844 Oustide_End:74455844 chro:chr2 SVtype:2 sup:2 Avg_Span:543 sumProb:2.000002
Inside_Start:106805021 Inside_End:106805021 OutSide_Start:107280900 Oustide_End:107280900 chro:chr14 SVtype:2 sup:2 Avg_Span:475879 sumProb:2.000002
Inside_Start:106809733 Inside_End:106809931 OutSide_Start:106810341 Oustide_End:106810366 chro:chr14 SVtype:2 sup:2 Avg_Span:521 sumProb:2.000002
Inside_Start:107169966 Inside_End:107169981 OutSide_Start:107170381 Oustide_End:107170418 chro:chr14 SVtype:2 sup:2 Avg_Span:426 sumProb:2.000001
Inside_Start:36048601 Inside_End:36048601 OutSide_Start:36049105 Oustide_End:36049105 chro:chr20 SVtype:2 sup:2 Avg_Span:504 sumProb:2.000001
Inside_Start:107065830 Inside_End:107065893 OutSide_Start:107066255 Oustide_End:107066327 chro:chr14 SVtype:2 sup:2 Avg_Span:429 sumProb:2.000000
Inside_Start:1278814 Inside_End:1278887 OutSide_Start:1279251 Oustide_End:1279352 chro:chr5 SVtype:2 sup:2 Avg_Span:451 sumProb:2.000000
Inside_Start:106572562 Inside_End:106572670 OutSide_Start:106573016 Oustide_End:106573074 chro:chr14 SVtype:2 sup:2 Avg_Span:429 sumProb:2.000000
TOTAL 6555
