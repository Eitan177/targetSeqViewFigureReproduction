HERE
1958
JJ
HH
Inside_Start:106518109 Inside_End:106518254 OutSide_Start:106573066 Oustide_End:106573254 chro:chr14 SVtype:2 sup:14 Avg_Span:54906 sumProb:inf
Inside_Start:106518116 Inside_End:106518240 OutSide_Start:107183212 Oustide_End:107183275 chro:chr14 SVtype:2 sup:10 Avg_Span:665042 sumProb:inf
Inside_Start:106626929 Inside_End:106627063 OutSide_Start:107074651 Oustide_End:107074791 chro:chr14 SVtype:2 sup:3 Avg_Span:447724 sumProb:inf
Inside_Start:106785365 Inside_End:106785586 OutSide_Start:106810129 Oustide_End:106810537 chro:chr14 SVtype:2 sup:5 Avg_Span:24776 sumProb:inf
Inside_Start:106805112 Inside_End:106805230 OutSide_Start:106877520 Oustide_End:106877655 chro:chr14 SVtype:2 sup:42 Avg_Span:72418 sumProb:inf
Inside_Start:106805010 Inside_End:106805228 OutSide_Start:107083049 Oustide_End:107083402 chro:chr14 SVtype:2 sup:18 Avg_Span:278095 sumProb:inf
Inside_Start:106823015 Inside_End:106823093 OutSide_Start:107273672 Oustide_End:107273732 chro:chr14 SVtype:2 sup:8 Avg_Span:450658 sumProb:inf
Inside_Start:106866319 Inside_End:106866363 OutSide_Start:107130925 Oustide_End:107131033 chro:chr14 SVtype:2 sup:8 Avg_Span:264598 sumProb:inf
Inside_Start:106993692 Inside_End:106993773 OutSide_Start:107183258 Oustide_End:107183298 chro:chr14 SVtype:2 sup:5 Avg_Span:189530 sumProb:inf
Inside_Start:22465891 Inside_End:22466108 OutSide_Start:22482793 Oustide_End:22482977 chro:chr15 SVtype:2 sup:6 Avg_Span:16890 sumProb:inf
Inside_Start:32859089 Inside_End:32859672 OutSide_Start:33815661 Oustide_End:33815731 chro:chr16 SVtype:4 sup:10 Avg_Span:956161 sumProb:inf
Inside_Start:32909563 Inside_End:32909566 OutSide_Start:33764079 Oustide_End:33764091 chro:chr16 SVtype:5 sup:2 Avg_Span:854520 sumProb:inf
Inside_Start:89442080 Inside_End:89442081 OutSide_Start:90078289 Oustide_End:90078289 chro:chr2 SVtype:4 sup:3 Avg_Span:636208 sumProb:inf
Inside_Start:89520749 Inside_End:89521145 OutSide_Start:89999416 Oustide_End:89999598 chro:chr2 SVtype:4 sup:3 Avg_Span:478605 sumProb:inf
Inside_Start:89513144 Inside_End:89513221 OutSide_Start:90249356 Oustide_End:90249420 chro:chr2 SVtype:5 sup:6 Avg_Span:736208 sumProb:inf
Inside_Start:107087099 Inside_End:107087212 OutSide_Start:107099109 Oustide_End:107099371 chro:chr14 SVtype:2 sup:19 Avg_Span:12006 sumProb:16.926514
Inside_Start:89161181 Inside_End:89161358 OutSide_Start:89901802 Oustide_End:89901927 chro:chr2 SVtype:5 sup:24 Avg_Span:740637 sumProb:15.452045
Inside_Start:106691357 Inside_End:106691549 OutSide_Start:107183249 Oustide_End:107183275 chro:chr14 SVtype:2 sup:6 Avg_Span:491766 sumProb:6.000000
Inside_Start:32993847 Inside_End:32994202 OutSide_Start:33673405 Oustide_End:33673773 chro:chr16 SVtype:4 sup:8 Avg_Span:679667 sumProb:4.446763
Inside_Start:33630287 Inside_End:33630287 OutSide_Start:33647227 Oustide_End:33647228 chro:chr16 SVtype:5 sup:4 Avg_Span:16940 sumProb:3.995469
Inside_Start:110547513 Inside_End:110547513 OutSide_Start:111339132 Oustide_End:111339132 chro:chr2 SVtype:4 sup:4 Avg_Span:791619 sumProb:3.831538
Inside_Start:33021059 Inside_End:33021120 OutSide_Start:33647074 Oustide_End:33647133 chro:chr16 SVtype:4 sup:9 Avg_Span:626023 sumProb:3.374441
Inside_Start:22298196 Inside_End:22298196 OutSide_Start:22555223 Oustide_End:22555223 chro:chr14 SVtype:2 sup:3 Avg_Span:257027 sumProb:3.000000
Inside_Start:1278342 Inside_End:1278449 OutSide_Start:1278786 Oustide_End:1278892 chro:chr5 SVtype:2 sup:3 Avg_Span:430 sumProb:3.000000
Inside_Start:142139104 Inside_End:142139273 OutSide_Start:142157325 Oustide_End:142157381 chro:chr7 SVtype:2 sup:3 Avg_Span:18183 sumProb:3.000000
Inside_Start:89495624 Inside_End:89495638 OutSide_Start:89986901 Oustide_End:89986969 chro:chr2 SVtype:4 sup:3 Avg_Span:491290 sumProb:2.997721
Inside_Start:89265663 Inside_End:89265800 OutSide_Start:89345426 Oustide_End:89345579 chro:chr2 SVtype:2 sup:4 Avg_Span:79775 sumProb:2.996626
Inside_Start:107094870 Inside_End:107095061 OutSide_Start:107280870 Oustide_End:107280893 chro:chr14 SVtype:2 sup:7 Avg_Span:185899 sumProb:2.545049
Inside_Start:106823028 Inside_End:106823042 OutSide_Start:107106296 Oustide_End:107106538 chro:chr14 SVtype:2 sup:3 Avg_Span:283360 sumProb:2.000796
Inside_Start:106559380 Inside_End:106559527 OutSide_Start:107178975 Oustide_End:107179107 chro:chr14 SVtype:2 sup:2 Avg_Span:619587 sumProb:2.000367
TOTAL 517
