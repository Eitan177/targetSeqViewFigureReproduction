HERE
1826
JJ
HH
Inside_Start:106466372 Inside_End:106466948 OutSide_Start:106466950 Oustide_End:106467755 chro:chr14 SVtype:2 sup:19 Avg_Span:635 sumProb:inf
Inside_Start:106518198 Inside_End:106518392 OutSide_Start:106993635 Oustide_End:106993946 chro:chr14 SVtype:2 sup:12 Avg_Span:475517 sumProb:inf
Inside_Start:106691357 Inside_End:106691668 OutSide_Start:106993616 Oustide_End:106993896 chro:chr14 SVtype:2 sup:5 Avg_Span:302254 sumProb:inf
Inside_Start:106785338 Inside_End:106785663 OutSide_Start:106810118 Oustide_End:106810560 chro:chr14 SVtype:2 sup:14 Avg_Span:24821 sumProb:inf
Inside_Start:106993601 Inside_End:106993724 OutSide_Start:107183199 Oustide_End:107183341 chro:chr14 SVtype:2 sup:16 Avg_Span:189564 sumProb:inf
Inside_Start:107048375 Inside_End:107048608 OutSide_Start:107130903 Oustide_End:107130959 chro:chr14 SVtype:2 sup:21 Avg_Span:82418 sumProb:inf
Inside_Start:32909241 Inside_End:32909271 OutSide_Start:33764190 Oustide_End:33764222 chro:chr16 SVtype:4 sup:7 Avg_Span:854936 sumProb:inf
Inside_Start:32993986 Inside_End:32994492 OutSide_Start:33673372 Oustide_End:33673771 chro:chr16 SVtype:4 sup:5 Avg_Span:679437 sumProb:inf
Inside_Start:32926961 Inside_End:32926972 OutSide_Start:33740685 Oustide_End:33740701 chro:chr16 SVtype:5 sup:7 Avg_Span:813731 sumProb:inf
Inside_Start:89521086 Inside_End:89521204 OutSide_Start:89999537 Oustide_End:89999652 chro:chr2 SVtype:4 sup:5 Avg_Span:478472 sumProb:inf
Inside_Start:142099503 Inside_End:142099503 OutSide_Start:142247274 Oustide_End:142247276 chro:chr7 SVtype:2 sup:2 Avg_Span:147772 sumProb:inf
Inside_Start:142131350 Inside_End:142131354 OutSide_Start:142148883 Oustide_End:142148899 chro:chr7 SVtype:2 sup:2 Avg_Span:17539 sumProb:inf
Inside_Start:142148958 Inside_End:142148981 OutSide_Start:142242456 Oustide_End:142242464 chro:chr7 SVtype:2 sup:2 Avg_Span:93490 sumProb:inf
Inside_Start:106691330 Inside_End:106691656 OutSide_Start:107183244 Oustide_End:107183280 chro:chr14 SVtype:2 sup:31 Avg_Span:491785 sumProb:29.984131
Inside_Start:107087136 Inside_End:107087324 OutSide_Start:107099206 Oustide_End:107099446 chro:chr14 SVtype:2 sup:15 Avg_Span:12069 sumProb:13.496533
Inside_Start:89161542 Inside_End:89161625 OutSide_Start:89185688 Oustide_End:89185835 chro:chr2 SVtype:5 sup:12 Avg_Span:24164 sumProb:12.000000
Inside_Start:107078149 Inside_End:107078379 OutSide_Start:107083255 Oustide_End:107083434 chro:chr14 SVtype:2 sup:21 Avg_Span:5011 sumProb:11.997589
Inside_Start:106559379 Inside_End:106559528 OutSide_Start:107178785 Oustide_End:107178989 chro:chr14 SVtype:2 sup:9 Avg_Span:619370 sumProb:9.000710
Inside_Start:106478112 Inside_End:106478145 OutSide_Start:106877659 Oustide_End:106877705 chro:chr14 SVtype:2 sup:10 Avg_Span:399548 sumProb:8.999605
Inside_Start:106330337 Inside_End:106330460 OutSide_Start:106354416 Oustide_End:106354668 chro:chr14 SVtype:2 sup:8 Avg_Span:24069 sumProb:8.000000
Inside_Start:106572839 Inside_End:106572948 OutSide_Start:107183194 Oustide_End:107183309 chro:chr14 SVtype:2 sup:10 Avg_Span:610355 sumProb:7.945440
Inside_Start:89533456 Inside_End:89533653 OutSide_Start:89976262 Oustide_End:89976399 chro:chr2 SVtype:4 sup:24 Avg_Span:442781 sumProb:7.691933
Inside_Start:23029810 Inside_End:23029873 OutSide_Start:23090492 Oustide_End:23090758 chro:chr22 SVtype:2 sup:6 Avg_Span:60805 sumProb:5.999966
Inside_Start:106477950 Inside_End:106478085 OutSide_Start:106829605 Oustide_End:106829673 chro:chr14 SVtype:2 sup:7 Avg_Span:351617 sumProb:5.969475
Inside_Start:106823022 Inside_End:106823047 OutSide_Start:107106289 Oustide_End:107106476 chro:chr14 SVtype:2 sup:6 Avg_Span:283358 sumProb:3.458660
Inside_Start:106466484 Inside_End:106466489 OutSide_Start:106467564 Oustide_End:106467703 chro:chr14 SVtype:2 sup:3 Avg_Span:1124 sumProb:3.024862
Inside_Start:106538996 Inside_End:106538996 OutSide_Start:107159851 Oustide_End:107159851 chro:chr14 SVtype:2 sup:3 Avg_Span:620855 sumProb:3.000000
Inside_Start:142099433 Inside_End:142099433 OutSide_Start:142119787 Oustide_End:142119787 chro:chr7 SVtype:2 sup:3 Avg_Span:20354 sumProb:3.000000
Inside_Start:106329376 Inside_End:106329413 OutSide_Start:106351893 Oustide_End:106351951 chro:chr14 SVtype:2 sup:3 Avg_Span:22511 sumProb:2.998802
Inside_Start:89512779 Inside_End:89512882 OutSide_Start:90007758 Oustide_End:90008286 chro:chr2 SVtype:4 sup:10 Avg_Span:495380 sumProb:2.584802
Inside_Start:89475624 Inside_End:89475782 OutSide_Start:89999344 Oustide_End:89999442 chro:chr2 SVtype:4 sup:7 Avg_Span:523671 sumProb:2.403609
Inside_Start:106804956 Inside_End:106805218 OutSide_Start:107083248 Oustide_End:107083273 chro:chr14 SVtype:2 sup:12 Avg_Span:278103 sumProb:2.070942
TOTAL 501
