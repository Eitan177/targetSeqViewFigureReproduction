HERE
1553
JJ
HH
Inside_Start:42385708 Inside_End:42385727 OutSide_Start:42387004 Oustide_End:42387433 chro:chr10 SVtype:2 sup:3 Avg_Span:1432 sumProb:inf
Inside_Start:42387770 Inside_End:42387780 OutSide_Start:42389494 Oustide_End:42389498 chro:chr10 SVtype:2 sup:3 Avg_Span:1722 sumProb:inf
Inside_Start:106691330 Inside_End:106691667 OutSide_Start:107183124 Oustide_End:107183291 chro:chr14 SVtype:2 sup:23 Avg_Span:491793 sumProb:inf
Inside_Start:106785330 Inside_End:106785421 OutSide_Start:106810119 Oustide_End:106810151 chro:chr14 SVtype:2 sup:16 Avg_Span:24738 sumProb:inf
Inside_Start:107078136 Inside_End:107078384 OutSide_Start:107083247 Oustide_End:107083407 chro:chr14 SVtype:2 sup:27 Avg_Span:4993 sumProb:inf
Inside_Start:32859603 Inside_End:32859673 OutSide_Start:33815661 Oustide_End:33815730 chro:chr16 SVtype:4 sup:10 Avg_Span:956072 sumProb:inf
Inside_Start:32990286 Inside_End:32990440 OutSide_Start:33677280 Oustide_End:33677939 chro:chr16 SVtype:5 sup:2 Avg_Span:687246 sumProb:inf
Inside_Start:107087147 Inside_End:107087262 OutSide_Start:107099203 Oustide_End:107099432 chro:chr14 SVtype:2 sup:4 Avg_Span:12110 sumProb:3.998715
Inside_Start:106798499 Inside_End:106798540 OutSide_Start:106823158 Oustide_End:106823697 chro:chr14 SVtype:2 sup:11 Avg_Span:24671 sumProb:2.501902
Inside_Start:23241267 Inside_End:23241770 OutSide_Start:23246946 Oustide_End:23247039 chro:chr22 SVtype:2 sup:4 Avg_Span:5411 sumProb:2.093937
Inside_Start:106933777 Inside_End:106933778 OutSide_Start:107175390 Oustide_End:107175469 chro:chr14 SVtype:2 sup:2 Avg_Span:241652 sumProb:2.033004
Inside_Start:106993732 Inside_End:106993732 OutSide_Start:107183280 Oustide_End:107183280 chro:chr14 SVtype:2 sup:2 Avg_Span:189548 sumProb:2.000011
TOTAL 245
