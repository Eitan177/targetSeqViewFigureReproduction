HERE
2984
JJ
HH
Inside_Start:122899739 Inside_End:122899739 OutSide_Start:123214985 Oustide_End:123214985 chro:chr11 SVtype:2 sup:2 Avg_Span:315246 sumProb:inf
Inside_Start:106466208 Inside_End:106466761 OutSide_Start:106466924 Oustide_End:106467800 chro:chr14 SVtype:2 sup:14 Avg_Span:721 sumProb:inf
Inside_Start:106466488 Inside_End:106466952 OutSide_Start:106467507 Oustide_End:106467734 chro:chr14 SVtype:2 sup:34 Avg_Span:675 sumProb:inf
Inside_Start:106466736 Inside_End:106466736 OutSide_Start:107147560 Oustide_End:107147560 chro:chr14 SVtype:2 sup:1 Avg_Span:680824 sumProb:inf
Inside_Start:106477967 Inside_End:106478176 OutSide_Start:106829616 Oustide_End:106829691 chro:chr14 SVtype:2 sup:35 Avg_Span:351576 sumProb:inf
Inside_Start:106518145 Inside_End:106518248 OutSide_Start:106691565 Oustide_End:106691699 chro:chr14 SVtype:2 sup:11 Avg_Span:173391 sumProb:inf
Inside_Start:106518049 Inside_End:106518246 OutSide_Start:106993594 Oustide_End:106993898 chro:chr14 SVtype:2 sup:8 Avg_Span:475507 sumProb:inf
Inside_Start:106552178 Inside_End:106552289 OutSide_Start:106926089 Oustide_End:106926257 chro:chr14 SVtype:2 sup:2 Avg_Span:373939 sumProb:inf
Inside_Start:106572919 Inside_End:106572947 OutSide_Start:107183219 Oustide_End:107183237 chro:chr14 SVtype:2 sup:3 Avg_Span:610296 sumProb:inf
Inside_Start:106626918 Inside_End:106627057 OutSide_Start:107074692 Oustide_End:107074778 chro:chr14 SVtype:2 sup:4 Avg_Span:447777 sumProb:inf
Inside_Start:106785238 Inside_End:106785612 OutSide_Start:106810118 Oustide_End:106810543 chro:chr14 SVtype:2 sup:16 Avg_Span:24756 sumProb:inf
Inside_Start:106805050 Inside_End:106805180 OutSide_Start:106877535 Oustide_End:106877659 chro:chr14 SVtype:2 sup:24 Avg_Span:72441 sumProb:inf
Inside_Start:106866156 Inside_End:106866392 OutSide_Start:107048526 Oustide_End:107048723 chro:chr14 SVtype:2 sup:18 Avg_Span:182285 sumProb:inf
Inside_Start:106993686 Inside_End:106993720 OutSide_Start:107183252 Oustide_End:107183596 chro:chr14 SVtype:2 sup:15 Avg_Span:189597 sumProb:inf
Inside_Start:107087224 Inside_End:107087247 OutSide_Start:107113939 Oustide_End:107114006 chro:chr14 SVtype:2 sup:3 Avg_Span:26741 sumProb:inf
Inside_Start:107106274 Inside_End:107106454 OutSide_Start:107273670 Oustide_End:107273700 chro:chr14 SVtype:2 sup:6 Avg_Span:167296 sumProb:inf
Inside_Start:32859126 Inside_End:32859651 OutSide_Start:33815603 Oustide_End:33815731 chro:chr16 SVtype:4 sup:11 Avg_Span:956175 sumProb:inf
Inside_Start:33630332 Inside_End:33630339 OutSide_Start:33661322 Oustide_End:33661386 chro:chr16 SVtype:5 sup:3 Avg_Span:31009 sumProb:inf
Inside_Start:89442110 Inside_End:89442110 OutSide_Start:90078262 Oustide_End:90078262 chro:chr2 SVtype:4 sup:5 Avg_Span:636152 sumProb:inf
Inside_Start:89521194 Inside_End:89521240 OutSide_Start:89999501 Oustide_End:89999543 chro:chr2 SVtype:4 sup:2 Avg_Span:478305 sumProb:inf
Inside_Start:89596915 Inside_End:89597173 OutSide_Start:89923871 Oustide_End:89924134 chro:chr2 SVtype:4 sup:3 Avg_Span:327044 sumProb:inf
Inside_Start:38374534 Inside_End:38374619 OutSide_Start:38380128 Oustide_End:38380444 chro:chr7 SVtype:2 sup:2 Avg_Span:5709 sumProb:inf
Inside_Start:106691330 Inside_End:106691555 OutSide_Start:107183226 Oustide_End:107183280 chro:chr14 SVtype:2 sup:38 Avg_Span:491791 sumProb:38.000004
Inside_Start:23029810 Inside_End:23029871 OutSide_Start:23090509 Oustide_End:23090737 chro:chr22 SVtype:2 sup:7 Avg_Span:60779 sumProb:6.999990
Inside_Start:106877360 Inside_End:106877637 OutSide_Start:107083051 Oustide_End:107083276 chro:chr14 SVtype:2 sup:19 Avg_Span:205711 sumProb:5.158515
Inside_Start:107239207 Inside_End:107239210 OutSide_Start:107239739 Oustide_End:107239921 chro:chr14 SVtype:2 sup:5 Avg_Span:605 sumProb:5.000000
Inside_Start:106653183 Inside_End:106653391 OutSide_Start:106845287 Oustide_End:106845409 chro:chr14 SVtype:2 sup:6 Avg_Span:192024 sumProb:4.998762
Inside_Start:107048562 Inside_End:107048637 OutSide_Start:107130949 Oustide_End:107131027 chro:chr14 SVtype:2 sup:5 Avg_Span:82393 sumProb:4.289477
Inside_Start:106559377 Inside_End:106559528 OutSide_Start:107178846 Oustide_End:107179093 chro:chr14 SVtype:2 sup:4 Avg_Span:619419 sumProb:4.000000
Inside_Start:22465960 Inside_End:22466012 OutSide_Start:22482835 Oustide_End:22482899 chro:chr15 SVtype:2 sup:4 Avg_Span:16865 sumProb:4.000000
Inside_Start:106798408 Inside_End:106798540 OutSide_Start:106823158 Oustide_End:106823616 chro:chr14 SVtype:2 sup:14 Avg_Span:24692 sumProb:3.003880
Inside_Start:142139141 Inside_End:142139141 OutSide_Start:142157207 Oustide_End:142157207 chro:chr7 SVtype:2 sup:3 Avg_Span:18066 sumProb:3.000032
Inside_Start:106478115 Inside_End:106478169 OutSide_Start:106877683 Oustide_End:106877707 chro:chr14 SVtype:2 sup:3 Avg_Span:399546 sumProb:3.000030
Inside_Start:106518038 Inside_End:106518330 OutSide_Start:106573064 Oustide_End:106573171 chro:chr14 SVtype:2 sup:8 Avg_Span:54921 sumProb:3.000003
Inside_Start:89533713 Inside_End:89533713 OutSide_Start:90091888 Oustide_End:90091888 chro:chr2 SVtype:4 sup:3 Avg_Span:558175 sumProb:2.999999
Inside_Start:106674801 Inside_End:106674801 OutSide_Start:107048549 Oustide_End:107048550 chro:chr14 SVtype:2 sup:3 Avg_Span:373748 sumProb:2.997718
Inside_Start:106805015 Inside_End:106805202 OutSide_Start:107083050 Oustide_End:107083356 chro:chr14 SVtype:2 sup:14 Avg_Span:278134 sumProb:2.834208
Inside_Start:106798290 Inside_End:106798312 OutSide_Start:107106281 Oustide_End:107106477 chro:chr14 SVtype:2 sup:5 Avg_Span:308028 sumProb:2.500001
Inside_Start:106691366 Inside_End:106691663 OutSide_Start:106993614 Oustide_End:106993898 chro:chr14 SVtype:2 sup:6 Avg_Span:302238 sumProb:2.000124
Inside_Start:142111151 Inside_End:142111280 OutSide_Start:142148792 Oustide_End:142148829 chro:chr7 SVtype:2 sup:2 Avg_Span:37595 sumProb:2.000124
Inside_Start:106780258 Inside_End:106780321 OutSide_Start:107095041 Oustide_End:107095046 chro:chr14 SVtype:2 sup:3 Avg_Span:314744 sumProb:2.000002
Inside_Start:23055690 Inside_End:23055753 OutSide_Start:23115042 Oustide_End:23115130 chro:chr22 SVtype:2 sup:3 Avg_Span:59389 sumProb:2.000001
TOTAL 709
