HERE
3391
JJ
HH
Inside_Start:106466393 Inside_End:106466968 OutSide_Start:106467211 Oustide_End:106467865 chro:chr14 SVtype:2 sup:30 Avg_Span:683 sumProb:inf
Inside_Start:106477939 Inside_End:106478176 OutSide_Start:106829607 Oustide_End:106829671 chro:chr14 SVtype:2 sup:31 Avg_Span:351582 sumProb:inf
Inside_Start:106477965 Inside_End:106478145 OutSide_Start:106780308 Oustide_End:106780785 chro:chr14 SVtype:2 sup:29 Avg_Span:302449 sumProb:inf
Inside_Start:106477992 Inside_End:106478118 OutSide_Start:106804992 Oustide_End:106805201 chro:chr14 SVtype:2 sup:6 Avg_Span:327017 sumProb:inf
Inside_Start:106518152 Inside_End:106518491 OutSide_Start:107183202 Oustide_End:107183656 chro:chr14 SVtype:2 sup:70 Avg_Span:665070 sumProb:inf
Inside_Start:106626895 Inside_End:106627056 OutSide_Start:107074647 Oustide_End:107074845 chro:chr14 SVtype:2 sup:9 Avg_Span:447749 sumProb:inf
Inside_Start:106691271 Inside_End:106691603 OutSide_Start:107183244 Oustide_End:107183458 chro:chr14 SVtype:2 sup:73 Avg_Span:491808 sumProb:inf
Inside_Start:106691278 Inside_End:106691674 OutSide_Start:106993606 Oustide_End:106993860 chro:chr14 SVtype:2 sup:11 Avg_Span:302266 sumProb:inf
Inside_Start:106780434 Inside_End:106780434 OutSide_Start:106877537 Oustide_End:106877612 chro:chr14 SVtype:2 sup:4 Avg_Span:97135 sumProb:inf
Inside_Start:106785336 Inside_End:106785421 OutSide_Start:106810117 Oustide_End:106810526 chro:chr14 SVtype:2 sup:25 Avg_Span:24748 sumProb:inf
Inside_Start:106798297 Inside_End:106798329 OutSide_Start:107106306 Oustide_End:107106549 chro:chr14 SVtype:2 sup:10 Avg_Span:308077 sumProb:inf
Inside_Start:106823004 Inside_End:106823229 OutSide_Start:107273627 Oustide_End:107273702 chro:chr14 SVtype:2 sup:3 Avg_Span:450541 sumProb:inf
Inside_Start:106993681 Inside_End:106993731 OutSide_Start:107183248 Oustide_End:107183303 chro:chr14 SVtype:2 sup:10 Avg_Span:189579 sumProb:inf
Inside_Start:107136523 Inside_End:107136540 OutSide_Start:107159792 Oustide_End:107159912 chro:chr14 SVtype:2 sup:2 Avg_Span:23320 sumProb:inf
Inside_Start:32926934 Inside_End:32927016 OutSide_Start:33740646 Oustide_End:33740727 chro:chr16 SVtype:5 sup:11 Avg_Span:813700 sumProb:inf
Inside_Start:23063398 Inside_End:23063619 OutSide_Start:23241801 Oustide_End:23242073 chro:chr22 SVtype:2 sup:6 Avg_Span:178383 sumProb:inf
Inside_Start:142099474 Inside_End:142099500 OutSide_Start:142247273 Oustide_End:142247305 chro:chr7 SVtype:2 sup:3 Avg_Span:147798 sumProb:inf
Inside_Start:142111063 Inside_End:142111350 OutSide_Start:142148822 Oustide_End:142148870 chro:chr7 SVtype:2 sup:4 Avg_Span:37605 sumProb:inf
Inside_Start:106330290 Inside_End:106330478 OutSide_Start:106357567 Oustide_End:106357746 chro:chr14 SVtype:2 sup:29 Avg_Span:27226 sumProb:29.000000
Inside_Start:106572840 Inside_End:106573093 OutSide_Start:107183211 Oustide_End:107183329 chro:chr14 SVtype:2 sup:14 Avg_Span:610351 sumProb:12.000085
Inside_Start:106372606 Inside_End:106372806 OutSide_Start:106382455 Oustide_End:106382623 chro:chr14 SVtype:2 sup:10 Avg_Span:9757 sumProb:9.972753
Inside_Start:1278294 Inside_End:1278569 OutSide_Start:1278729 Oustide_End:1279001 chro:chr5 SVtype:2 sup:8 Avg_Span:451 sumProb:8.000000
Inside_Start:22465921 Inside_End:22466103 OutSide_Start:22482813 Oustide_End:22483271 chro:chr15 SVtype:2 sup:10 Avg_Span:16956 sumProb:7.963373
Inside_Start:107087145 Inside_End:107087255 OutSide_Start:107099289 Oustide_End:107099386 chro:chr14 SVtype:2 sup:9 Avg_Span:12120 sumProb:7.003222
Inside_Start:106466237 Inside_End:106466761 OutSide_Start:106467274 Oustide_End:106467891 chro:chr14 SVtype:2 sup:9 Avg_Span:1068 sumProb:6.480261
Inside_Start:106470872 Inside_End:106471123 OutSide_Start:107078212 Oustide_End:107078343 chro:chr14 SVtype:2 sup:6 Avg_Span:607255 sumProb:6.000000
Inside_Start:106804944 Inside_End:106805306 OutSide_Start:107083034 Oustide_End:107083428 chro:chr14 SVtype:2 sup:26 Avg_Span:278145 sumProb:5.989269
Inside_Start:22298127 Inside_End:22298256 OutSide_Start:22418896 Oustide_End:22418959 chro:chr14 SVtype:2 sup:5 Avg_Span:120714 sumProb:5.000000
Inside_Start:106877372 Inside_End:106877649 OutSide_Start:107083200 Oustide_End:107083360 chro:chr14 SVtype:2 sup:14 Avg_Span:205692 sumProb:4.363831
Inside_Start:106798475 Inside_End:106798671 OutSide_Start:106798909 Oustide_End:106799100 chro:chr14 SVtype:2 sup:6 Avg_Span:448 sumProb:4.238414
Inside_Start:106467640 Inside_End:106467640 OutSide_Start:107218725 Oustide_End:107218725 chro:chr14 SVtype:2 sup:4 Avg_Span:751085 sumProb:4.000000
Inside_Start:106966808 Inside_End:106967039 OutSide_Start:106967216 Oustide_End:106967467 chro:chr14 SVtype:2 sup:4 Avg_Span:419 sumProb:4.000000
Inside_Start:106559527 Inside_End:106559528 OutSide_Start:107178829 Oustide_End:107179051 chro:chr14 SVtype:2 sup:4 Avg_Span:619392 sumProb:3.999992
Inside_Start:22461585 Inside_End:22461936 OutSide_Start:22462147 Oustide_End:22462438 chro:chr15 SVtype:2 sup:4 Avg_Span:495 sumProb:3.999798
Inside_Start:106787192 Inside_End:106787315 OutSide_Start:107022031 Oustide_End:107022123 chro:chr14 SVtype:2 sup:4 Avg_Span:234815 sumProb:3.996593
Inside_Start:89416657 Inside_End:89416715 OutSide_Start:90193282 Oustide_End:90193428 chro:chr2 SVtype:4 sup:5 Avg_Span:776722 sumProb:3.994673
Inside_Start:33020568 Inside_End:33021107 OutSide_Start:33647086 Oustide_End:33647121 chro:chr16 SVtype:4 sup:6 Avg_Span:626084 sumProb:3.621629
Inside_Start:107094852 Inside_End:107095022 OutSide_Start:107280871 Oustide_End:107280895 chro:chr14 SVtype:2 sup:11 Avg_Span:185938 sumProb:3.312048
Inside_Start:142143340 Inside_End:142143569 OutSide_Start:142180396 Oustide_End:142180428 chro:chr7 SVtype:2 sup:3 Avg_Span:36923 sumProb:3.026378
Inside_Start:106471071 Inside_End:106471100 OutSide_Start:107159727 Oustide_End:107159773 chro:chr14 SVtype:2 sup:3 Avg_Span:688652 sumProb:3.000000
Inside_Start:22294063 Inside_End:22294125 OutSide_Start:22294470 Oustide_End:22294557 chro:chr14 SVtype:2 sup:3 Avg_Span:429 sumProb:3.000000
Inside_Start:22977960 Inside_End:22978003 OutSide_Start:22978405 Oustide_End:22978452 chro:chr14 SVtype:2 sup:3 Avg_Span:446 sumProb:3.000000
Inside_Start:106620246 Inside_End:106620246 OutSide_Start:107055828 Oustide_End:107055828 chro:chr14 SVtype:2 sup:3 Avg_Span:435582 sumProb:3.000000
Inside_Start:106630740 Inside_End:106630791 OutSide_Start:107159890 Oustide_End:107159932 chro:chr14 SVtype:2 sup:3 Avg_Span:529161 sumProb:3.000000
Inside_Start:106773749 Inside_End:106773804 OutSide_Start:106774204 Oustide_End:106774209 chro:chr14 SVtype:2 sup:3 Avg_Span:431 sumProb:3.000000
Inside_Start:107078191 Inside_End:107078293 OutSide_Start:107159790 Oustide_End:107159946 chro:chr14 SVtype:2 sup:3 Avg_Span:81635 sumProb:3.000000
Inside_Start:107273479 Inside_End:107273789 OutSide_Start:107273943 Oustide_End:107274304 chro:chr14 SVtype:2 sup:3 Avg_Span:483 sumProb:3.000000
Inside_Start:38369708 Inside_End:38370009 OutSide_Start:38407260 Oustide_End:38407423 chro:chr7 SVtype:2 sup:3 Avg_Span:37460 sumProb:3.000000
Inside_Start:106578787 Inside_End:106578787 OutSide_Start:107078156 Oustide_End:107078157 chro:chr14 SVtype:2 sup:3 Avg_Span:499369 sumProb:2.999999
Inside_Start:23029820 Inside_End:23029869 OutSide_Start:23090528 Oustide_End:23090912 chro:chr22 SVtype:2 sup:4 Avg_Span:60879 sumProb:2.999993
Inside_Start:22265873 Inside_End:22266003 OutSide_Start:22372720 Oustide_End:22372822 chro:chr14 SVtype:2 sup:3 Avg_Span:106828 sumProb:2.999743
Inside_Start:106597943 Inside_End:106597943 OutSide_Start:106626967 Oustide_End:106626967 chro:chr14 SVtype:2 sup:3 Avg_Span:29024 sumProb:2.996626
Inside_Start:32050605 Inside_End:32050605 OutSide_Start:32916998 Oustide_End:32916998 chro:chr16 SVtype:2 sup:3 Avg_Span:866393 sumProb:2.996052
Inside_Start:107057135 Inside_End:107057254 OutSide_Start:107275805 Oustide_End:107275888 chro:chr14 SVtype:2 sup:3 Avg_Span:218672 sumProb:2.789606
Inside_Start:20210663 Inside_End:20211028 OutSide_Start:20211070 Oustide_End:20211449 chro:chr15 SVtype:2 sup:7 Avg_Span:425 sumProb:2.249343
Inside_Start:106962661 Inside_End:106962965 OutSide_Start:107169883 Oustide_End:107169983 chro:chr14 SVtype:2 sup:3 Avg_Span:207086 sumProb:2.147230
Inside_Start:89160650 Inside_End:89160756 OutSide_Start:89890899 Oustide_End:89891166 chro:chr2 SVtype:4 sup:4 Avg_Span:730307 sumProb:2.026357
Inside_Start:106493874 Inside_End:106494121 OutSide_Start:107178671 Oustide_End:107178934 chro:chr14 SVtype:2 sup:2 Avg_Span:684805 sumProb:2.006140
Inside_Start:106780282 Inside_End:106780348 OutSide_Start:106805107 Oustide_End:106805133 chro:chr14 SVtype:2 sup:4 Avg_Span:24801 sumProb:2.002293
Inside_Start:106471230 Inside_End:106471248 OutSide_Start:106539172 Oustide_End:106539296 chro:chr14 SVtype:2 sup:3 Avg_Span:67971 sumProb:2.001394
Inside_Start:106471178 Inside_End:106471229 OutSide_Start:107113789 Oustide_End:107113868 chro:chr14 SVtype:2 sup:2 Avg_Span:642625 sumProb:2.001078
Inside_Start:38369813 Inside_End:38369990 OutSide_Start:38402531 Oustide_End:38402610 chro:chr7 SVtype:2 sup:4 Avg_Span:32650 sumProb:2.000003
Inside_Start:106805015 Inside_End:106805111 OutSide_Start:107280846 Oustide_End:107280951 chro:chr14 SVtype:2 sup:3 Avg_Span:475853 sumProb:2.000000
TOTAL 1104
